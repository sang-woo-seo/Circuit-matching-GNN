.SUBCKT level_shift3 IN OUT VDD VBIASH VBIASL VSS
M1 tn1 tn2 VDD VDD PMOS W=3.5u L=350.00n M=1
M2 tn2 tn1 VDD VDD PMOS W=3.5u L=350.00n M=1
M3 tn3 VBIASH tn1 VDD PMOS W=3.5u L=350.00n M=1
M4 OUT VBIASH tn2 VDD PMOS W=3.5u L=350.00n M=1
M5 tn3 VBIASL tn5 VSS NMOS W=1.4u L=350.00n M=1
M6 OUT VBIASL tn6 VSS NMOS W=1.4u L=350.00n M=1
M7 tn5 INB VSS VSS NMOS W=1.4u L=350.00n M=1
M8 tn6 IN VSS VSS NMOS W=1.4u L=350.00n M=1
XIV1 IN INB inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
.ENDS
