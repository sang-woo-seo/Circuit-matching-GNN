.SUBCKT col_sel3_8m a<2> a<1> a<0> cs<7> cs<6> cs<5> cs<4> cs<3> cs<2> cs<1>
+cs<0> ena pre xvld
XI51 net33 net31 net25 ena pre cs<7> xvld   col_sel1m
XI41 net35 net29 net27 ena pre cs<0> xvld   col_sel1m
XI49 net35 net31 net27 ena pre cs<2> xvld   col_sel1m
XI50 net35 net31 net25 ena pre cs<6> xvld   col_sel1m
XI47 net33 net29 net27 ena pre cs<1> xvld   col_sel1m
XI52 net33 net29 net25 ena pre cs<5> xvld   col_sel1m
XI48 net33 net31 net27 ena pre cs<3> xvld   col_sel1m
XI53 net35 net29 net25 ena pre cs<4> xvld   col_sel1m
XI88 net35 net33   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI56 a<2> net27   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI90 a<0> net35   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI57 net27 net25   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI54 net29 net31   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI55 a<1> net29   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
.ENDS
