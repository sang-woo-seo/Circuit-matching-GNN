.SUBCKT ctrl256kbm a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8>
+a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> cs<511> cs<510> cs<509> cs<508>
+cs<507> cs<506> cs<505> cs<504> cs<503> cs<502> cs<501> cs<500> cs<499>
+cs<498> cs<497> cs<496> cs<495> cs<494> cs<493> cs<492> cs<491> cs<490>
+cs<489> cs<488> cs<487> cs<486> cs<485> cs<484> cs<483> cs<482> cs<481>
+cs<480> cs<479> cs<478> cs<477> cs<476> cs<475> cs<474> cs<473> cs<472>
+cs<471> cs<470> cs<469> cs<468> cs<467> cs<466> cs<465> cs<464> cs<463>
+cs<462> cs<461> cs<460> cs<459> cs<458> cs<457> cs<456> cs<455> cs<454>
+cs<453> cs<452> cs<451> cs<450> cs<449> cs<448> cs<447> cs<446> cs<445>
+cs<444> cs<443> cs<442> cs<441> cs<440> cs<439> cs<438> cs<437> cs<436>
+cs<435> cs<434> cs<433> cs<432> cs<431> cs<430> cs<429> cs<428> cs<427>
+cs<426> cs<425> cs<424> cs<423> cs<422> cs<421> cs<420> cs<419> cs<418>
+cs<417> cs<416> cs<415> cs<414> cs<413> cs<412> cs<411> cs<410> cs<409>
+cs<408> cs<407> cs<406> cs<405> cs<404> cs<403> cs<402> cs<401> cs<400>
+cs<399> cs<398> cs<397> cs<396> cs<395> cs<394> cs<393> cs<392> cs<391>
+cs<390> cs<389> cs<388> cs<387> cs<386> cs<385> cs<384> cs<383> cs<382>
+cs<381> cs<380> cs<379> cs<378> cs<377> cs<376> cs<375> cs<374> cs<373>
+cs<372> cs<371> cs<370> cs<369> cs<368> cs<367> cs<366> cs<365> cs<364>
+cs<363> cs<362> cs<361> cs<360> cs<359> cs<358> cs<357> cs<356> cs<355>
+cs<354> cs<353> cs<352> cs<351> cs<350> cs<349> cs<348> cs<347> cs<346>
+cs<345> cs<344> cs<343> cs<342> cs<341> cs<340> cs<339> cs<338> cs<337>
+cs<336> cs<335> cs<334> cs<333> cs<332> cs<331> cs<330> cs<329> cs<328>
+cs<327> cs<326> cs<325> cs<324> cs<323> cs<322> cs<321> cs<320> cs<319>
+cs<318> cs<317> cs<316> cs<315> cs<314> cs<313> cs<312> cs<311> cs<310>
+cs<309> cs<308> cs<307> cs<306> cs<305> cs<304> cs<303> cs<302> cs<301>
+cs<300> cs<299> cs<298> cs<297> cs<296> cs<295> cs<294> cs<293> cs<292>
+cs<291> cs<290> cs<289> cs<288> cs<287> cs<286> cs<285> cs<284> cs<283>
+cs<282> cs<281> cs<280> cs<279> cs<278> cs<277> cs<276> cs<275> cs<274>
+cs<273> cs<272> cs<271> cs<270> cs<269> cs<268> cs<267> cs<266> cs<265>
+cs<264> cs<263> cs<262> cs<261> cs<260> cs<259> cs<258> cs<257> cs<256>
+cs<255> cs<254> cs<253> cs<252> cs<251> cs<250> cs<249> cs<248> cs<247>
+cs<246> cs<245> cs<244> cs<243> cs<242> cs<241> cs<240> cs<239> cs<238>
+cs<237> cs<236> cs<235> cs<234> cs<233> cs<232> cs<231> cs<230> cs<229>
+cs<228> cs<227> cs<226> cs<225> cs<224> cs<223> cs<222> cs<221> cs<220>
+cs<219> cs<218> cs<217> cs<216> cs<215> cs<214> cs<213> cs<212> cs<211>
+cs<210> cs<209> cs<208> cs<207> cs<206> cs<205> cs<204> cs<203> cs<202>
+cs<201> cs<200> cs<199> cs<198> cs<197> cs<196> cs<195> cs<194> cs<193>
+cs<192> cs<191> cs<190> cs<189> cs<188> cs<187> cs<186> cs<185> cs<184>
+cs<183> cs<182> cs<181> cs<180> cs<179> cs<178> cs<177> cs<176> cs<175>
+cs<174> cs<173> cs<172> cs<171> cs<170> cs<169> cs<168> cs<167> cs<166>
+cs<165> cs<164> cs<163> cs<162> cs<161> cs<160> cs<159> cs<158> cs<157>
+cs<156> cs<155> cs<154> cs<153> cs<152> cs<151> cs<150> cs<149> cs<148>
+cs<147> cs<146> cs<145> cs<144> cs<143> cs<142> cs<141> cs<140> cs<139>
+cs<138> cs<137> cs<136> cs<135> cs<134> cs<133> cs<132> cs<131> cs<130>
+cs<129> cs<128> cs<127> cs<126> cs<125> cs<124> cs<123> cs<122> cs<121>
+cs<120> cs<119> cs<118> cs<117> cs<116> cs<115> cs<114> cs<113> cs<112>
+cs<111> cs<110> cs<109> cs<108> cs<107> cs<106> cs<105> cs<104> cs<103>
+cs<102> cs<101> cs<100> cs<99> cs<98> cs<97> cs<96> cs<95> cs<94> cs<93>
+cs<92> cs<91> cs<90> cs<89> cs<88> cs<87> cs<86> cs<85> cs<84> cs<83> cs<82>
+cs<81> cs<80> cs<79> cs<78> cs<77> cs<76> cs<75> cs<74> cs<73> cs<72> cs<71>
+cs<70> cs<69> cs<68> cs<67> cs<66> cs<65> cs<64> cs<63> cs<62> cs<61> cs<60>
+cs<59> cs<58> cs<57> cs<56> cs<55> cs<54> cs<53> cs<52> cs<51> cs<50> cs<49>
+cs<48> cs<47> cs<46> cs<45> cs<44> cs<43> cs<42> cs<41> cs<40> cs<39> cs<38>
+cs<37> cs<36> cs<35> cs<34> cs<33> cs<32> cs<31> cs<30> cs<29> cs<28> cs<27>
+cs<26> cs<25> cs<24> cs<23> cs<22> cs<21> cs<20> cs<19> cs<18> cs<17> cs<16>
+cs<15> cs<14> cs<13> cs<12> cs<11> cs<10> cs<9> cs<8> cs<7> cs<6> cs<5> cs<4>
+cs<3> cs<2> cs<1> cs<0> ena l_sel main_ena n_ena p_ena pre r_sel w_ wl<511>
+wl<510> wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502>
+wl<501> wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493>
+wl<492> wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484>
+wl<483> wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475>
+wl<474> wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466>
+wl<465> wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457>
+wl<456> wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448>
+wl<447> wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439>
+wl<438> wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430>
+wl<429> wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421>
+wl<420> wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412>
+wl<411> wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403>
+wl<402> wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394>
+wl<393> wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385>
+wl<384> wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376>
+wl<375> wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367>
+wl<366> wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358>
+wl<357> wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349>
+wl<348> wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340>
+wl<339> wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331>
+wl<330> wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322>
+wl<321> wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313>
+wl<312> wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304>
+wl<303> wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295>
+wl<294> wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286>
+wl<285> wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277>
+wl<276> wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268>
+wl<267> wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259>
+wl<258> wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250>
+wl<249> wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241>
+wl<240> wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232>
+wl<231> wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223>
+wl<222> wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214>
+wl<213> wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205>
+wl<204> wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196>
+wl<195> wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187>
+wl<186> wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178>
+wl<177> wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169>
+wl<168> wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160>
+wl<159> wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151>
+wl<150> wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142>
+wl<141> wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133>
+wl<132> wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124>
+wl<123> wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115>
+wl<114> wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106>
+wl<105> wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96>
+wl<95> wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85>
+wl<84> wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74>
+wl<73> wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63>
+wl<62> wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52>
+wl<51> wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41>
+wl<40> wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30>
+wl<29> wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19>
+wl<18> wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8>
+wl<7> wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>
XI139 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> ena w_ net107   atd18m
XI88 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> cs<511> cs<510>
+cs<509> cs<508> cs<507> cs<506> cs<505> cs<504> cs<503> cs<502> cs<501>
+cs<500> cs<499> cs<498> cs<497> cs<496> cs<495> cs<494> cs<493> cs<492>
+cs<491> cs<490> cs<489> cs<488> cs<487> cs<486> cs<485> cs<484> cs<483>
+cs<482> cs<481> cs<480> cs<479> cs<478> cs<477> cs<476> cs<475> cs<474>
+cs<473> cs<472> cs<471> cs<470> cs<469> cs<468> cs<467> cs<466> cs<465>
+cs<464> cs<463> cs<462> cs<461> cs<460> cs<459> cs<458> cs<457> cs<456>
+cs<455> cs<454> cs<453> cs<452> cs<451> cs<450> cs<449> cs<448> cs<447>
+cs<446> cs<445> cs<444> cs<443> cs<442> cs<441> cs<440> cs<439> cs<438>
+cs<437> cs<436> cs<435> cs<434> cs<433> cs<432> cs<431> cs<430> cs<429>
+cs<428> cs<427> cs<426> cs<425> cs<424> cs<423> cs<422> cs<421> cs<420>
+cs<419> cs<418> cs<417> cs<416> cs<415> cs<414> cs<413> cs<412> cs<411>
+cs<410> cs<409> cs<408> cs<407> cs<406> cs<405> cs<404> cs<403> cs<402>
+cs<401> cs<400> cs<399> cs<398> cs<397> cs<396> cs<395> cs<394> cs<393>
+cs<392> cs<391> cs<390> cs<389> cs<388> cs<387> cs<386> cs<385> cs<384>
+cs<383> cs<382> cs<381> cs<380> cs<379> cs<378> cs<377> cs<376> cs<375>
+cs<374> cs<373> cs<372> cs<371> cs<370> cs<369> cs<368> cs<367> cs<366>
+cs<365> cs<364> cs<363> cs<362> cs<361> cs<360> cs<359> cs<358> cs<357>
+cs<356> cs<355> cs<354> cs<353> cs<352> cs<351> cs<350> cs<349> cs<348>
+cs<347> cs<346> cs<345> cs<344> cs<343> cs<342> cs<341> cs<340> cs<339>
+cs<338> cs<337> cs<336> cs<335> cs<334> cs<333> cs<332> cs<331> cs<330>
+cs<329> cs<328> cs<327> cs<326> cs<325> cs<324> cs<323> cs<322> cs<321>
+cs<320> cs<319> cs<318> cs<317> cs<316> cs<315> cs<314> cs<313> cs<312>
+cs<311> cs<310> cs<309> cs<308> cs<307> cs<306> cs<305> cs<304> cs<303>
+cs<302> cs<301> cs<300> cs<299> cs<298> cs<297> cs<296> cs<295> cs<294>
+cs<293> cs<292> cs<291> cs<290> cs<289> cs<288> cs<287> cs<286> cs<285>
+cs<284> cs<283> cs<282> cs<281> cs<280> cs<279> cs<278> cs<277> cs<276>
+cs<275> cs<274> cs<273> cs<272> cs<271> cs<270> cs<269> cs<268> cs<267>
+cs<266> cs<265> cs<264> cs<263> cs<262> cs<261> cs<260> cs<259> cs<258>
+cs<257> cs<256> cs<255> cs<254> cs<253> cs<252> cs<251> cs<250> cs<249>
+cs<248> cs<247> cs<246> cs<245> cs<244> cs<243> cs<242> cs<241> cs<240>
+cs<239> cs<238> cs<237> cs<236> cs<235> cs<234> cs<233> cs<232> cs<231>
+cs<230> cs<229> cs<228> cs<227> cs<226> cs<225> cs<224> cs<223> cs<222>
+cs<221> cs<220> cs<219> cs<218> cs<217> cs<216> cs<215> cs<214> cs<213>
+cs<212> cs<211> cs<210> cs<209> cs<208> cs<207> cs<206> cs<205> cs<204>
+cs<203> cs<202> cs<201> cs<200> cs<199> cs<198> cs<197> cs<196> cs<195>
+cs<194> cs<193> cs<192> cs<191> cs<190> cs<189> cs<188> cs<187> cs<186>
+cs<185> cs<184> cs<183> cs<182> cs<181> cs<180> cs<179> cs<178> cs<177>
+cs<176> cs<175> cs<174> cs<173> cs<172> cs<171> cs<170> cs<169> cs<168>
+cs<167> cs<166> cs<165> cs<164> cs<163> cs<162> cs<161> cs<160> cs<159>
+cs<158> cs<157> cs<156> cs<155> cs<154> cs<153> cs<152> cs<151> cs<150>
+cs<149> cs<148> cs<147> cs<146> cs<145> cs<144> cs<143> cs<142> cs<141>
+cs<140> cs<139> cs<138> cs<137> cs<136> cs<135> cs<134> cs<133> cs<132>
+cs<131> cs<130> cs<129> cs<128> cs<127> cs<126> cs<125> cs<124> cs<123>
+cs<122> cs<121> cs<120> cs<119> cs<118> cs<117> cs<116> cs<115> cs<114>
+cs<113> cs<112> cs<111> cs<110> cs<109> cs<108> cs<107> cs<106> cs<105>
+cs<104> cs<103> cs<102> cs<101> cs<100> cs<99> cs<98> cs<97> cs<96> cs<95>
+cs<94> cs<93> cs<92> cs<91> cs<90> cs<89> cs<88> cs<87> cs<86> cs<85> cs<84>
+cs<83> cs<82> cs<81> cs<80> cs<79> cs<78> cs<77> cs<76> cs<75> cs<74> cs<73>
+cs<72> cs<71> cs<70> cs<69> cs<68> cs<67> cs<66> cs<65> cs<64> cs<63> cs<62>
+cs<61> cs<60> cs<59> cs<58> cs<57> cs<56> cs<55> cs<54> cs<53> cs<52> cs<51>
+cs<50> cs<49> cs<48> cs<47> cs<46> cs<45> cs<44> cs<43> cs<42> cs<41> cs<40>
+cs<39> cs<38> cs<37> cs<36> cs<35> cs<34> cs<33> cs<32> cs<31> cs<30> cs<29>
+cs<28> cs<27> cs<26> cs<25> cs<24> cs<23> cs<22> cs<21> cs<20> cs<19> cs<18>
+cs<17> cs<16> cs<15> cs<14> cs<13> cs<12> cs<11> cs<10> cs<9> cs<8> cs<7>
+cs<6> cs<5> cs<4> cs<3> cs<2> cs<1> cs<0> ena pre net102   col_sel9_512
XI58 a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> ena net107 wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0> xvld   deco9_512
XI99 net102 net75   delay4
XI97 xvld net77 net106 w_   ctg Lp=0.35u Wp=1.4u Ln=0.35u Wn=1.4u
XI96 net85 net77 w_ net106   ctg Lp=0.35u Wp=1.4u Ln=0.35u Wn=1.4u
XI90 xvld net85   delay10
XI146 net116 pre r_sel xvld   rl_sel
XI145 a<8> pre l_sel xvld   rl_sel
XI82 n_ena p_ena xvld   sen_ena
XI100 net75 net98   inv Ln=0.35u Wn=3.5u M=1 Lp=0.35u Wp=7u
XI101 net98 main_ena   inv Ln=0.35u Wn=3.5u M=3 Lp=0.35u Wp=7u
XI95 net104 net102   inv Ln=0.35u Wn=3.5u M=3 Lp=0.35u Wp=7u
XI94 net77 net104   inv Ln=0.35u Wn=3.5u M=1 Lp=0.35u Wp=7u
XI98 w_ net106   inv Ln=0.35u Wn=3.5u M=1 Lp=0.35u Wp=7u
XI108 net107 net108   inv Ln=0.35u Wn=36u M=2 Lp=0.35u Wp=72u
XI81 net114 xvld   inv Ln=0.35u Wn=10u M=9 Lp=0.35u Wp=20u
XI110 net108 pre   inv Ln=0.35u Wn=36u M=5 Lp=0.35u Wp=72u
XI80 net113 net114   inv Ln=0.35u Wn=10u M=3 Lp=0.35u Wp=20u
XI147 a<8> net116   inv Ln=0.35u Wn=3.5u M=1 Lp=0.35u Wp=7u
XI79 pre net113   xvald
.ENDS
