.SUBCKT level_shift2 IN OUT VDD VSS
M1 tn1 OUT VDD VDD PMOS W=3.5u L=350.00n M=1
M2 tn2 tn3 VDD VDD PMOS W=3.5u L=350.00n M=1
M3 tn3 IN tn1 VDD PMOS W=3.5u L=350.00n M=1
M4 OUT INB tn2 VDD PMOS W=3.5u L=350.00n M=1
M5 tn3 IN VSS VSS NMOS W=1.4u L=350.00n M=1
M6 OUT INB VSS VSS NMOS W=1.4u L=350.00n M=1
XIV1 IN INB inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
.ENDS
