.SUBCKT level_shift1 IN OUT VDD VSS
M1 tn1 OUT VDD VDD PMOS W=3.5u L=350.00n M=1
M2 OUT tn1 VDD VDD PMOS W=3.5u L=350.00n M=1
M3 tn1 IN VSS VSS NMOS W=1.4u L=350.00n M=1
M4 OUT INB VSS VSS NMOS W=1.4u L=350.00n M=1
XIV1 IN INB inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
.ENDS
