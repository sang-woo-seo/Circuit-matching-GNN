.SUBCKT sa_pre bl blb br brb cs io io_ l_sel n_ena p_ena pre r_sel
MM11 net51 net40 net039 vdd! PMOS W=14u L=350.00n M=1
MM15 net40 net51 net039 vdd! PMOS W=14u L=350.00n M=1
MM12 vdd! p_ena net039 vdd! PMOS W=14u L=350.00n M=1
MM80 bl pre blb vbb! NMOS W=1.4u L=350.00n M=1
MM81 vddh! pre blb vbb! NMOS W=1.4u L=350.00n M=1
MM82 vddh! pre bl vbb! NMOS W=1.4u L=350.00n M=1
MM73 br pre brb vbb! NMOS W=1.4u L=350.00n M=1
MM72 vddh! pre br vbb! NMOS W=1.4u L=350.00n M=1
MM71 vddh! pre brb vbb! NMOS W=1.4u L=350.00n M=1
MM76 net40 pre net51 vbb! NMOS W=1.4u L=350.00n M=1
MM75 vddh! pre net40 vbb! NMOS W=1.4u L=350.00n M=1
MM0 blb l_sel net51 vbb! NMOS W=1.4u L=350.00n M=1
MM1 bl l_sel net40 vbb! NMOS W=1.4u L=350.00n M=1
MM77 net51 net40 net081 vbb! NMOS W=7u L=350.00n M=1
MM78 net081 n_ena gnd! vbb! NMOS W=7u L=350.00n M=1
MM79 net40 net51 net081 vbb! NMOS W=7u L=350.00n M=1
MM7 net40 r_sel br vbb! NMOS W=1.4u L=350.00n M=1
MM8 net51 r_sel brb vbb! NMOS W=1.4u L=350.00n M=1
MM9 net40 cs io vbb! NMOS W=1.4u L=350.00n M=1
MM10 io_ cs net51 vbb! NMOS W=1.4u L=350.00n M=1
MM74 vddh! pre net51 vbb! NMOS W=1.4u L=350.00n M=1
.ENDS
