.SUBCKT col_sel9_512 a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> cs<511>
+cs<510> cs<509> cs<508> cs<507> cs<506> cs<505> cs<504> cs<503> cs<502>
+cs<501> cs<500> cs<499> cs<498> cs<497> cs<496> cs<495> cs<494> cs<493>
+cs<492> cs<491> cs<490> cs<489> cs<488> cs<487> cs<486> cs<485> cs<484>
+cs<483> cs<482> cs<481> cs<480> cs<479> cs<478> cs<477> cs<476> cs<475>
+cs<474> cs<473> cs<472> cs<471> cs<470> cs<469> cs<468> cs<467> cs<466>
+cs<465> cs<464> cs<463> cs<462> cs<461> cs<460> cs<459> cs<458> cs<457>
+cs<456> cs<455> cs<454> cs<453> cs<452> cs<451> cs<450> cs<449> cs<448>
+cs<447> cs<446> cs<445> cs<444> cs<443> cs<442> cs<441> cs<440> cs<439>
+cs<438> cs<437> cs<436> cs<435> cs<434> cs<433> cs<432> cs<431> cs<430>
+cs<429> cs<428> cs<427> cs<426> cs<425> cs<424> cs<423> cs<422> cs<421>
+cs<420> cs<419> cs<418> cs<417> cs<416> cs<415> cs<414> cs<413> cs<412>
+cs<411> cs<410> cs<409> cs<408> cs<407> cs<406> cs<405> cs<404> cs<403>
+cs<402> cs<401> cs<400> cs<399> cs<398> cs<397> cs<396> cs<395> cs<394>
+cs<393> cs<392> cs<391> cs<390> cs<389> cs<388> cs<387> cs<386> cs<385>
+cs<384> cs<383> cs<382> cs<381> cs<380> cs<379> cs<378> cs<377> cs<376>
+cs<375> cs<374> cs<373> cs<372> cs<371> cs<370> cs<369> cs<368> cs<367>
+cs<366> cs<365> cs<364> cs<363> cs<362> cs<361> cs<360> cs<359> cs<358>
+cs<357> cs<356> cs<355> cs<354> cs<353> cs<352> cs<351> cs<350> cs<349>
+cs<348> cs<347> cs<346> cs<345> cs<344> cs<343> cs<342> cs<341> cs<340>
+cs<339> cs<338> cs<337> cs<336> cs<335> cs<334> cs<333> cs<332> cs<331>
+cs<330> cs<329> cs<328> cs<327> cs<326> cs<325> cs<324> cs<323> cs<322>
+cs<321> cs<320> cs<319> cs<318> cs<317> cs<316> cs<315> cs<314> cs<313>
+cs<312> cs<311> cs<310> cs<309> cs<308> cs<307> cs<306> cs<305> cs<304>
+cs<303> cs<302> cs<301> cs<300> cs<299> cs<298> cs<297> cs<296> cs<295>
+cs<294> cs<293> cs<292> cs<291> cs<290> cs<289> cs<288> cs<287> cs<286>
+cs<285> cs<284> cs<283> cs<282> cs<281> cs<280> cs<279> cs<278> cs<277>
+cs<276> cs<275> cs<274> cs<273> cs<272> cs<271> cs<270> cs<269> cs<268>
+cs<267> cs<266> cs<265> cs<264> cs<263> cs<262> cs<261> cs<260> cs<259>
+cs<258> cs<257> cs<256> cs<255> cs<254> cs<253> cs<252> cs<251> cs<250>
+cs<249> cs<248> cs<247> cs<246> cs<245> cs<244> cs<243> cs<242> cs<241>
+cs<240> cs<239> cs<238> cs<237> cs<236> cs<235> cs<234> cs<233> cs<232>
+cs<231> cs<230> cs<229> cs<228> cs<227> cs<226> cs<225> cs<224> cs<223>
+cs<222> cs<221> cs<220> cs<219> cs<218> cs<217> cs<216> cs<215> cs<214>
+cs<213> cs<212> cs<211> cs<210> cs<209> cs<208> cs<207> cs<206> cs<205>
+cs<204> cs<203> cs<202> cs<201> cs<200> cs<199> cs<198> cs<197> cs<196>
+cs<195> cs<194> cs<193> cs<192> cs<191> cs<190> cs<189> cs<188> cs<187>
+cs<186> cs<185> cs<184> cs<183> cs<182> cs<181> cs<180> cs<179> cs<178>
+cs<177> cs<176> cs<175> cs<174> cs<173> cs<172> cs<171> cs<170> cs<169>
+cs<168> cs<167> cs<166> cs<165> cs<164> cs<163> cs<162> cs<161> cs<160>
+cs<159> cs<158> cs<157> cs<156> cs<155> cs<154> cs<153> cs<152> cs<151>
+cs<150> cs<149> cs<148> cs<147> cs<146> cs<145> cs<144> cs<143> cs<142>
+cs<141> cs<140> cs<139> cs<138> cs<137> cs<136> cs<135> cs<134> cs<133>
+cs<132> cs<131> cs<130> cs<129> cs<128> cs<127> cs<126> cs<125> cs<124>
+cs<123> cs<122> cs<121> cs<120> cs<119> cs<118> cs<117> cs<116> cs<115>
+cs<114> cs<113> cs<112> cs<111> cs<110> cs<109> cs<108> cs<107> cs<106>
+cs<105> cs<104> cs<103> cs<102> cs<101> cs<100> cs<99> cs<98> cs<97> cs<96>
+cs<95> cs<94> cs<93> cs<92> cs<91> cs<90> cs<89> cs<88> cs<87> cs<86> cs<85>
+cs<84> cs<83> cs<82> cs<81> cs<80> cs<79> cs<78> cs<77> cs<76> cs<75> cs<74>
+cs<73> cs<72> cs<71> cs<70> cs<69> cs<68> cs<67> cs<66> cs<65> cs<64> cs<63>
+cs<62> cs<61> cs<60> cs<59> cs<58> cs<57> cs<56> cs<55> cs<54> cs<53> cs<52>
+cs<51> cs<50> cs<49> cs<48> cs<47> cs<46> cs<45> cs<44> cs<43> cs<42> cs<41>
+cs<40> cs<39> cs<38> cs<37> cs<36> cs<35> cs<34> cs<33> cs<32> cs<31> cs<30>
+cs<29> cs<28> cs<27> cs<26> cs<25> cs<24> cs<23> cs<22> cs<21> cs<20> cs<19>
+cs<18> cs<17> cs<16> cs<15> cs<14> cs<13> cs<12> cs<11> cs<10> cs<9> cs<8>
+cs<7> cs<6> cs<5> cs<4> cs<3> cs<2> cs<1> cs<0> ena pre xvld
XI63 a<6> a<5> a<4> a<3> a<2> a<1> a<0> cs<127> cs<126> cs<125> cs<124>
+cs<123> cs<122> cs<121> cs<120> cs<119> cs<118> cs<117> cs<116> cs<115>
+cs<114> cs<113> cs<112> cs<111> cs<110> cs<109> cs<108> cs<107> cs<106>
+cs<105> cs<104> cs<103> cs<102> cs<101> cs<100> cs<99> cs<98> cs<97> cs<96>
+cs<95> cs<94> cs<93> cs<92> cs<91> cs<90> cs<89> cs<88> cs<87> cs<86> cs<85>
+cs<84> cs<83> cs<82> cs<81> cs<80> cs<79> cs<78> cs<77> cs<76> cs<75> cs<74>
+cs<73> cs<72> cs<71> cs<70> cs<69> cs<68> cs<67> cs<66> cs<65> cs<64> cs<63>
+cs<62> cs<61> cs<60> cs<59> cs<58> cs<57> cs<56> cs<55> cs<54> cs<53> cs<52>
+cs<51> cs<50> cs<49> cs<48> cs<47> cs<46> cs<45> cs<44> cs<43> cs<42> cs<41>
+cs<40> cs<39> cs<38> cs<37> cs<36> cs<35> cs<34> cs<33> cs<32> cs<31> cs<30>
+cs<29> cs<28> cs<27> cs<26> cs<25> cs<24> cs<23> cs<22> cs<21> cs<20> cs<19>
+cs<18> cs<17> cs<16> cs<15> cs<14> cs<13> cs<12> cs<11> cs<10> cs<9> cs<8>
+cs<7> cs<6> cs<5> cs<4> cs<3> cs<2> cs<1> cs<0> net<0> net110 net108  
+col_sel7_128
XI66 a<6> a<5> a<4> a<3> a<2> a<1> a<0> cs<511> cs<510> cs<509> cs<508>
+cs<507> cs<506> cs<505> cs<504> cs<503> cs<502> cs<501> cs<500> cs<499>
+cs<498> cs<497> cs<496> cs<495> cs<494> cs<493> cs<492> cs<491> cs<490>
+cs<489> cs<488> cs<487> cs<486> cs<485> cs<484> cs<483> cs<482> cs<481>
+cs<480> cs<479> cs<478> cs<477> cs<476> cs<475> cs<474> cs<473> cs<472>
+cs<471> cs<470> cs<469> cs<468> cs<467> cs<466> cs<465> cs<464> cs<463>
+cs<462> cs<461> cs<460> cs<459> cs<458> cs<457> cs<456> cs<455> cs<454>
+cs<453> cs<452> cs<451> cs<450> cs<449> cs<448> cs<447> cs<446> cs<445>
+cs<444> cs<443> cs<442> cs<441> cs<440> cs<439> cs<438> cs<437> cs<436>
+cs<435> cs<434> cs<433> cs<432> cs<431> cs<430> cs<429> cs<428> cs<427>
+cs<426> cs<425> cs<424> cs<423> cs<422> cs<421> cs<420> cs<419> cs<418>
+cs<417> cs<416> cs<415> cs<414> cs<413> cs<412> cs<411> cs<410> cs<409>
+cs<408> cs<407> cs<406> cs<405> cs<404> cs<403> cs<402> cs<401> cs<400>
+cs<399> cs<398> cs<397> cs<396> cs<395> cs<394> cs<393> cs<392> cs<391>
+cs<390> cs<389> cs<388> cs<387> cs<386> cs<385> cs<384> net<3> net110 net108
+  col_sel7_128
XI65 a<6> a<5> a<4> a<3> a<2> a<1> a<0> cs<383> cs<382> cs<381> cs<380>
+cs<379> cs<378> cs<377> cs<376> cs<375> cs<374> cs<373> cs<372> cs<371>
+cs<370> cs<369> cs<368> cs<367> cs<366> cs<365> cs<364> cs<363> cs<362>
+cs<361> cs<360> cs<359> cs<358> cs<357> cs<356> cs<355> cs<354> cs<353>
+cs<352> cs<351> cs<350> cs<349> cs<348> cs<347> cs<346> cs<345> cs<344>
+cs<343> cs<342> cs<341> cs<340> cs<339> cs<338> cs<337> cs<336> cs<335>
+cs<334> cs<333> cs<332> cs<331> cs<330> cs<329> cs<328> cs<327> cs<326>
+cs<325> cs<324> cs<323> cs<322> cs<321> cs<320> cs<319> cs<318> cs<317>
+cs<316> cs<315> cs<314> cs<313> cs<312> cs<311> cs<310> cs<309> cs<308>
+cs<307> cs<306> cs<305> cs<304> cs<303> cs<302> cs<301> cs<300> cs<299>
+cs<298> cs<297> cs<296> cs<295> cs<294> cs<293> cs<292> cs<291> cs<290>
+cs<289> cs<288> cs<287> cs<286> cs<285> cs<284> cs<283> cs<282> cs<281>
+cs<280> cs<279> cs<278> cs<277> cs<276> cs<275> cs<274> cs<273> cs<272>
+cs<271> cs<270> cs<269> cs<268> cs<267> cs<266> cs<265> cs<264> cs<263>
+cs<262> cs<261> cs<260> cs<259> cs<258> cs<257> cs<256> net<2> net110 net108
+  col_sel7_128
XI64 a<6> a<5> a<4> a<3> a<2> a<1> a<0> cs<255> cs<254> cs<253> cs<252>
+cs<251> cs<250> cs<249> cs<248> cs<247> cs<246> cs<245> cs<244> cs<243>
+cs<242> cs<241> cs<240> cs<239> cs<238> cs<237> cs<236> cs<235> cs<234>
+cs<233> cs<232> cs<231> cs<230> cs<229> cs<228> cs<227> cs<226> cs<225>
+cs<224> cs<223> cs<222> cs<221> cs<220> cs<219> cs<218> cs<217> cs<216>
+cs<215> cs<214> cs<213> cs<212> cs<211> cs<210> cs<209> cs<208> cs<207>
+cs<206> cs<205> cs<204> cs<203> cs<202> cs<201> cs<200> cs<199> cs<198>
+cs<197> cs<196> cs<195> cs<194> cs<193> cs<192> cs<191> cs<190> cs<189>
+cs<188> cs<187> cs<186> cs<185> cs<184> cs<183> cs<182> cs<181> cs<180>
+cs<179> cs<178> cs<177> cs<176> cs<175> cs<174> cs<173> cs<172> cs<171>
+cs<170> cs<169> cs<168> cs<167> cs<166> cs<165> cs<164> cs<163> cs<162>
+cs<161> cs<160> cs<159> cs<158> cs<157> cs<156> cs<155> cs<154> cs<153>
+cs<152> cs<151> cs<150> cs<149> cs<148> cs<147> cs<146> cs<145> cs<144>
+cs<143> cs<142> cs<141> cs<140> cs<139> cs<138> cs<137> cs<136> cs<135>
+cs<134> cs<133> cs<132> cs<131> cs<130> cs<129> cs<128> net<1> net110 net108
+  col_sel7_128
XI61 a<8> a<7> ena net<3> net<2> net<1> net<0>   decoder2_4
XI55 pre net112   inv Ln=0.35u Wn=8u M=9 Lp=0.35u Wp=16u
XI54 net112 net110   inv Ln=0.35u Wn=8u M=27 Lp=0.35u Wp=16u
XI79 net106 net108   inv Ln=0.35u Wn=8u M=6 Lp=0.35u Wp=16u
XI80 xvld net106   inv Ln=0.35u Wn=10u M=2 Lp=0.35u Wp=20u
.ENDS
