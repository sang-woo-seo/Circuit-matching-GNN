.SUBCKT main_sense ena io io_ o o_ pre
XI165 pre net20   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
MM5 o pre o_ vbb! NMOS W=1.4u L=350.00n M=1
MM2 o_ io net21 vbb! NMOS W=7u L=350.00n M=1
MM3 o io_ net21 vbb! NMOS W=7u L=350.00n M=1
MM4 net21 ena gnd! vbb! NMOS W=7u L=350.00n M=1
MM0 vdd! o_ o vdd! PMOS W=14u L=350.00n M=1
MM1 o_ net20 o vdd! PMOS W=1.4u L=350.00n M=1
MM17 vdd! o o_ vdd! PMOS W=14u L=350.00n M=1
.ENDS
