.SUBCKT deco9_512 a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> ena pre wl<511>
+wl<510> wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502>
+wl<501> wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493>
+wl<492> wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484>
+wl<483> wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475>
+wl<474> wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466>
+wl<465> wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457>
+wl<456> wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448>
+wl<447> wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439>
+wl<438> wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430>
+wl<429> wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421>
+wl<420> wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412>
+wl<411> wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403>
+wl<402> wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394>
+wl<393> wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385>
+wl<384> wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376>
+wl<375> wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367>
+wl<366> wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358>
+wl<357> wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349>
+wl<348> wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340>
+wl<339> wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331>
+wl<330> wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322>
+wl<321> wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313>
+wl<312> wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304>
+wl<303> wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295>
+wl<294> wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286>
+wl<285> wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277>
+wl<276> wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268>
+wl<267> wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259>
+wl<258> wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250>
+wl<249> wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241>
+wl<240> wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232>
+wl<231> wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223>
+wl<222> wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214>
+wl<213> wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205>
+wl<204> wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196>
+wl<195> wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187>
+wl<186> wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178>
+wl<177> wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169>
+wl<168> wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160>
+wl<159> wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151>
+wl<150> wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142>
+wl<141> wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133>
+wl<132> wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124>
+wl<123> wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115>
+wl<114> wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106>
+wl<105> wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96>
+wl<95> wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85>
+wl<84> wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74>
+wl<73> wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63>
+wl<62> wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52>
+wl<51> wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41>
+wl<40> wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30>
+wl<29> wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19>
+wl<18> wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8>
+wl<7> wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0> xvld
XI61 a<8> a<7> ena net<3> net<2> net<1> net<0>   decoder2_4
XI63 a<6> a<5> a<4> a<3> a<2> a<1> a<0> net<0> net110 wl<127> wl<126> wl<125>
+wl<124> wl<123> wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116>
+wl<115> wl<114> wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107>
+wl<106> wl<105> wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97>
+wl<96> wl<95> wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86>
+wl<85> wl<84> wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75>
+wl<74> wl<73> wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64>
+wl<63> wl<62> wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53>
+wl<52> wl<51> wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42>
+wl<41> wl<40> wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31>
+wl<30> wl<29> wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20>
+wl<19> wl<18> wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9>
+wl<8> wl<7> wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0> net108   deco7_128
XI66 a<6> a<5> a<4> a<3> a<2> a<1> a<0> net<3> net110 wl<511> wl<510> wl<509>
+wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501> wl<500>
+wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492> wl<491>
+wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483> wl<482>
+wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474> wl<473>
+wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465> wl<464>
+wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456> wl<455>
+wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447> wl<446>
+wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438> wl<437>
+wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429> wl<428>
+wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420> wl<419>
+wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411> wl<410>
+wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402> wl<401>
+wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393> wl<392>
+wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384> net108  
+deco7_128
XI65 a<6> a<5> a<4> a<3> a<2> a<1> a<0> net<2> net110 wl<383> wl<382> wl<381>
+wl<380> wl<379> wl<378> wl<377> wl<376> wl<375> wl<374> wl<373> wl<372>
+wl<371> wl<370> wl<369> wl<368> wl<367> wl<366> wl<365> wl<364> wl<363>
+wl<362> wl<361> wl<360> wl<359> wl<358> wl<357> wl<356> wl<355> wl<354>
+wl<353> wl<352> wl<351> wl<350> wl<349> wl<348> wl<347> wl<346> wl<345>
+wl<344> wl<343> wl<342> wl<341> wl<340> wl<339> wl<338> wl<337> wl<336>
+wl<335> wl<334> wl<333> wl<332> wl<331> wl<330> wl<329> wl<328> wl<327>
+wl<326> wl<325> wl<324> wl<323> wl<322> wl<321> wl<320> wl<319> wl<318>
+wl<317> wl<316> wl<315> wl<314> wl<313> wl<312> wl<311> wl<310> wl<309>
+wl<308> wl<307> wl<306> wl<305> wl<304> wl<303> wl<302> wl<301> wl<300>
+wl<299> wl<298> wl<297> wl<296> wl<295> wl<294> wl<293> wl<292> wl<291>
+wl<290> wl<289> wl<288> wl<287> wl<286> wl<285> wl<284> wl<283> wl<282>
+wl<281> wl<280> wl<279> wl<278> wl<277> wl<276> wl<275> wl<274> wl<273>
+wl<272> wl<271> wl<270> wl<269> wl<268> wl<267> wl<266> wl<265> wl<264>
+wl<263> wl<262> wl<261> wl<260> wl<259> wl<258> wl<257> wl<256> net108  
+deco7_128
XI64 a<6> a<5> a<4> a<3> a<2> a<1> a<0> net<1> net110 wl<255> wl<254> wl<253>
+wl<252> wl<251> wl<250> wl<249> wl<248> wl<247> wl<246> wl<245> wl<244>
+wl<243> wl<242> wl<241> wl<240> wl<239> wl<238> wl<237> wl<236> wl<235>
+wl<234> wl<233> wl<232> wl<231> wl<230> wl<229> wl<228> wl<227> wl<226>
+wl<225> wl<224> wl<223> wl<222> wl<221> wl<220> wl<219> wl<218> wl<217>
+wl<216> wl<215> wl<214> wl<213> wl<212> wl<211> wl<210> wl<209> wl<208>
+wl<207> wl<206> wl<205> wl<204> wl<203> wl<202> wl<201> wl<200> wl<199>
+wl<198> wl<197> wl<196> wl<195> wl<194> wl<193> wl<192> wl<191> wl<190>
+wl<189> wl<188> wl<187> wl<186> wl<185> wl<184> wl<183> wl<182> wl<181>
+wl<180> wl<179> wl<178> wl<177> wl<176> wl<175> wl<174> wl<173> wl<172>
+wl<171> wl<170> wl<169> wl<168> wl<167> wl<166> wl<165> wl<164> wl<163>
+wl<162> wl<161> wl<160> wl<159> wl<158> wl<157> wl<156> wl<155> wl<154>
+wl<153> wl<152> wl<151> wl<150> wl<149> wl<148> wl<147> wl<146> wl<145>
+wl<144> wl<143> wl<142> wl<141> wl<140> wl<139> wl<138> wl<137> wl<136>
+wl<135> wl<134> wl<133> wl<132> wl<131> wl<130> wl<129> wl<128> net108  
+deco7_128
XI55 pre net112   inv Ln=0.35u Wn=8u M=9 Lp=0.35u Wp=16u
XI54 net112 net110   inv Ln=0.35u Wn=8u M=27 Lp=0.35u Wp=16u
XI79 net106 net108   inv Ln=0.35u Wn=8u M=6 Lp=0.35u Wp=16u
XI80 xvld net106   inv Ln=0.35u Wn=10u M=2 Lp=0.35u Wp=20u
.ENDS
