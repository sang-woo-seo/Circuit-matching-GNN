.SUBCKT deco7_128 a<6> a<5> a<4> a<3> a<2> a<1> a<0> ena pre wl<127> wl<126>
+wl<125> wl<124> wl<123> wl<122> wl<121> wl<120> wl<119> wl<118> wl<117>
+wl<116> wl<115> wl<114> wl<113> wl<112> wl<111> wl<110> wl<109> wl<108>
+wl<107> wl<106> wl<105> wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98>
+wl<97> wl<96> wl<95> wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87>
+wl<86> wl<85> wl<84> wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76>
+wl<75> wl<74> wl<73> wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65>
+wl<64> wl<63> wl<62> wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54>
+wl<53> wl<52> wl<51> wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43>
+wl<42> wl<41> wl<40> wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32>
+wl<31> wl<30> wl<29> wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21>
+wl<20> wl<19> wl<18> wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10>
+wl<9> wl<8> wl<7> wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0> xvld
XI61 a<6> a<5> a<4> a<3> ena net<15> net<14> net<13> net<12> net<11> net<10>
+net<9> net<8> net<7> net<6> net<5> net<4> net<3> net<2> net<1> net<0>  
+decoder4_16
XI81 pre net199   inv Ln=0.35u Wn=8u M=27 Lp=0.35u Wp=16u
XI84 xvld net211   inv Ln=0.35u Wn=10u M=6 Lp=0.35u Wp=20u
XI55 pre net112   inv Ln=0.35u Wn=8u M=27 Lp=0.35u Wp=16u
XI54 net112 net110   inv Ln=0.35u Wn=8u M=81 Lp=0.35u Wp=16u
XI82 net199 net201   inv Ln=0.35u Wn=8u M=81 Lp=0.35u Wp=16u
XI79 net106 net108   inv Ln=0.35u Wn=10u M=18 Lp=0.35u Wp=20u
XI80 xvld net106   inv Ln=0.35u Wn=10u M=6 Lp=0.35u Wp=20u
XI83 net211 net213   inv Ln=0.35u Wn=10u M=18 Lp=0.35u Wp=20u
XI72 a<2> a<1> a<0> net<15> net201 wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> net213   deco3_8m
XI73 a<2> a<1> a<0> net<11> net201 wl<95> wl<94> wl<93> wl<92> wl<91> wl<90>
+wl<89> wl<88> net213   deco3_8m
XI74 a<2> a<1> a<0> net<10> net201 wl<87> wl<86> wl<85> wl<84> wl<83> wl<82>
+wl<81> wl<80> net213   deco3_8m
XI75 a<2> a<1> a<0> net<9> net201 wl<79> wl<78> wl<77> wl<76> wl<75> wl<74>
+wl<73> wl<72> net213   deco3_8m
XI76 a<2> a<1> a<0> net<12> net201 wl<103> wl<102> wl<101> wl<100> wl<99>
+wl<98> wl<97> wl<96> net213   deco3_8m
XI77 a<2> a<1> a<0> net<14> net201 wl<119> wl<118> wl<117> wl<116> wl<115>
+wl<114> wl<113> wl<112> net213   deco3_8m
XI78 a<2> a<1> a<0> net<13> net201 wl<111> wl<110> wl<109> wl<108> wl<107>
+wl<106> wl<105> wl<104> net213   deco3_8m
XI71 a<2> a<1> a<0> net<8> net201 wl<71> wl<70> wl<69> wl<68> wl<67> wl<66>
+wl<65> wl<64> net213   deco3_8m
XI63 a<2> a<1> a<0> net<0> net110 wl<7> wl<6> wl<5> wl<4> wl<3> wl<2> wl<1>
+wl<0> net108   deco3_8m
XI70 a<2> a<1> a<0> net<7> net110 wl<63> wl<62> wl<61> wl<60> wl<59> wl<58>
+wl<57> wl<56> net108   deco3_8m
XI66 a<2> a<1> a<0> net<3> net110 wl<31> wl<30> wl<29> wl<28> wl<27> wl<26>
+wl<25> wl<24> net108   deco3_8m
XI65 a<2> a<1> a<0> net<2> net110 wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> net108   deco3_8m
XI64 a<2> a<1> a<0> net<1> net110 wl<15> wl<14> wl<13> wl<12> wl<11> wl<10>
+wl<9> wl<8> net108   deco3_8m
XI67 a<2> a<1> a<0> net<4> net110 wl<39> wl<38> wl<37> wl<36> wl<35> wl<34>
+wl<33> wl<32> net108   deco3_8m
XI69 a<2> a<1> a<0> net<6> net110 wl<55> wl<54> wl<53> wl<52> wl<51> wl<50>
+wl<49> wl<48> net108   deco3_8m
XI68 a<2> a<1> a<0> net<5> net110 wl<47> wl<46> wl<45> wl<44> wl<43> wl<42>
+wl<41> wl<40> net108   deco3_8m
.ENDS
