.SUBCKT bank16mx1n a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14>
+a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> ena
+i_o w_
XI66 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<22> i_o w_   block512x512n
XI65 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<6> i_o w_   block512x512n
XI64 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<23> i_o w_   block512x512n
XI63 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<7> i_o w_   block512x512n
XI62 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<8> i_o w_   block512x512n
XI61 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<25> i_o w_   block512x512n
XI59 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<27> i_o w_   block512x512n
XI58 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<24> i_o w_   block512x512n
XI57 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<20> i_o w_   block512x512n
XI56 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<21> i_o w_   block512x512n
XI55 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<26> i_o w_   block512x512n
XI54 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<4> i_o w_   block512x512n
XI53 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<11> i_o w_   block512x512n
XI52 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<5> i_o w_   block512x512n
XI49 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<10> i_o w_   block512x512n
XI35 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<39> i_o w_   block512x512n
XI36 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<40> i_o w_   block512x512n
XI41 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<52> i_o w_   block512x512n
XI32 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<54> i_o w_   block512x512n
XI47 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<41> i_o w_   block512x512n
XI51 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<9> i_o w_   block512x512n
XI38 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<59> i_o w_   block512x512n
XI48 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<42> i_o w_   block512x512n
XI18 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<33> i_o w_   block512x512n
XI21 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<62> i_o w_   block512x512n
XI20 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<32> i_o w_   block512x512n
XI42 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<53> i_o w_   block512x512n
XI22 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<49> i_o w_   block512x512n
XI28 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<35> i_o w_   block512x512n
XI31 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<50> i_o w_   block512x512n
XI27 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<44> i_o w_   block512x512n
XI25 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<63> i_o w_   block512x512n
XI30 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<34> i_o w_   block512x512n
XI19 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<47> i_o w_   block512x512n
XI26 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<61> i_o w_   block512x512n
XI24 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<60> i_o w_   block512x512n
XI34 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<55> i_o w_   block512x512n
XI23 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<48> i_o w_   block512x512n
XI17 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<45> i_o w_   block512x512n
XI3 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<14> i_o w_   block512x512n
XI5 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<13> i_o w_   block512x512n
XI2 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<1> i_o w_   block512x512n
XI1 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<15> i_o w_   block512x512n
XI0 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<0> i_o w_   block512x512n
XI11 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<30> i_o w_   block512x512n
XI10 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<17> i_o w_   block512x512n
XI8 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<16> i_o w_   block512x512n
XI15 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<28> i_o w_   block512x512n
XI9 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<31> i_o w_   block512x512n
XI13 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<29> i_o w_   block512x512n
XI7 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<12> i_o w_   block512x512n
XI6 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<3> i_o w_   block512x512n
XI14 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<19> i_o w_   block512x512n
XI4 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<2> i_o w_   block512x512n
XI12 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<18> i_o w_   block512x512n
XI39 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<56> i_o w_   block512x512n
XI16 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<46> i_o w_   block512x512n
XI37 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<57> i_o w_   block512x512n
XI29 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<51> i_o w_   block512x512n
XI43 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<58> i_o w_   block512x512n
XI45 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<43> i_o w_   block512x512n
XI46 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<37> i_o w_   block512x512n
XI33 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<38> i_o w_   block512x512n
XI44 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<36> i_o w_   block512x512n
XI68 a<23> a<22> a<21> a<20> a<19> a<18> ena en<63> en<62> en<61> en<60>
+en<59> en<58> en<57> en<56> en<55> en<54> en<53> en<52> en<51> en<50> en<49>
+en<48> en<47> en<46> en<45> en<44> en<43> en<42> en<41> en<40> en<39> en<38>
+en<37> en<36> en<35> en<34> en<33> en<32> en<31> en<30> en<29> en<28> en<27>
+en<26> en<25> en<24> en<23> en<22> en<21> en<20> en<19> en<18> en<17> en<16>
+en<15> en<14> en<13> en<12> en<11> en<10> en<9> en<8> en<7> en<6> en<5> en<4>
+en<3> en<2> en<1> en<0>   decoder6_64
.ENDS
