.SUBCKT decoder6_64 A<5> A<4> A<3> A<2> A<1> A<0> ENA X<63> X<62> X<61> X<60>
+X<59> X<58> X<57> X<56> X<55> X<54> X<53> X<52> X<51> X<50> X<49> X<48> X<47>
+X<46> X<45> X<44> X<43> X<42> X<41> X<40> X<39> X<38> X<37> X<36> X<35> X<34>
+X<33> X<32> X<31> X<30> X<29> X<28> X<27> X<26> X<25> X<24> X<23> X<22> X<21>
+X<20> X<19> X<18> X<17> X<16> X<15> X<14> X<13> X<12> X<11> X<10> X<9> X<8>
+X<7> X<6> X<5> X<4> X<3> X<2> X<1> X<0>
XI95 A<5> A<4> ENA en<3> en<2> en<1> en<0>   decoder2_4
XI97 A<3> A<2> A<1> A<0> en<2> X<47> X<46> X<45> X<44> X<43> X<42> X<41> X<40>
+X<39> X<38> X<37> X<36> X<35> X<34> X<33> X<32>   decoder4_16
XI98 A<3> A<2> A<1> A<0> en<3> X<63> X<62> X<61> X<60> X<59> X<58> X<57> X<56>
+X<55> X<54> X<53> X<52> X<51> X<50> X<49> X<48>   decoder4_16
XI94 A<3> A<2> A<1> A<0> en<0> X<15> X<14> X<13> X<12> X<11> X<10> X<9> X<8>
+X<7> X<6> X<5> X<4> X<3> X<2> X<1> X<0>   decoder4_16
XI96 A<3> A<2> A<1> A<0> en<1> X<31> X<30> X<29> X<28> X<27> X<26> X<25> X<24>
+X<23> X<22> X<21> X<20> X<19> X<18> X<17> X<16>   decoder4_16
.ENDS
