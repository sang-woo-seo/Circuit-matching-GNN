.SUBCKT nand5 A B C D E Y
MM3 net40 D net12 vbb! NMOS W=Wn L=Ln M=1
MM1 net60 C net40 vbb! NMOS W=Wn L=Ln M=1
MM14 net28 B net60 vbb! NMOS W=Wn L=Ln M=1
MM13 Y A net28 vbb! NMOS W=Wn L=Ln M=1
MM4 net12 E gnd! vbb! NMOS W=Wn L=Ln M=1
MM5 Y E vdd! vdd! PMOS W=Wp L=Lp M=1
MM2 Y D vdd! vdd! PMOS W=Wp L=Lp M=1
MM0 Y C vdd! vdd! PMOS W=Wp L=Lp M=1
MM12 Y A vdd! vdd! PMOS W=Wp L=Lp M=1
MM11 Y B vdd! vdd! PMOS W=Wp L=Lp M=1
.ENDS
