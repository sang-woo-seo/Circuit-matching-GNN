.SUBCKT array512x1 cs io io_ l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>
XI817 bl vddh! wl<307>   mc
XI584 br vddh! wl<133>   mc
XI607 blb vddh! wl<388>   mc
XI813 bl vddh! wl<309>   mc
XI585 brb vddh! wl<128>   mc
XI662 blb vddh! wl<490>   mc
XI680 blb vddh! wl<508>   mc
XI579 br vddh! wl<129>   mc
XI636 bl vddh! wl<447>   mc
XI586 brb vddh! wl<130>   mc
XI639 blb vddh! wl<442>   mc
XI653 blb vddh! wl<428>   mc
XI763 bl vddh! wl<381>   mc
XI587 br vddh! wl<141>   mc
XI757 blb vddh! wl<374>   mc
XI488 brb vddh! wl<220>   mc
XI511 brb vddh! wl<250>   mc
XI582 brb vddh! wl<132>   mc
XI828 bl vddh! wl<287>   mc
XI519 br vddh! wl<231>   mc
XI588 br vddh! wl<143>   mc
XI741 bl vddh! wl<345>   mc
XI789 bl vddh! wl<297>   mc
XI559 brb vddh! wl<180>   mc
XI577 brb vddh! wl<152>   mc
XI578 br vddh! wl<155>   mc
XI567 br vddh! wl<151>   mc
XI589 brb vddh! wl<140>   mc
XI645 blb vddh! wl<422>   mc
XI838 blb vddh! wl<260>   mc
XI661 bl vddh! wl<489>   mc
XI580 br vddh! wl<131>   mc
XI850 bl vddh! wl<267>   mc
XI576 br vddh! wl<153>   mc
XI581 brb vddh! wl<134>   mc
XI583 br vddh! wl<135>   mc
XI575 brb vddh! wl<154>   mc
XI613 bl vddh! wl<409>   mc
XI748 blb vddh! wl<336>   mc
XI535 brb vddh! wl<174>   mc
XI753 bl vddh! wl<339>   mc
XI772 bl vddh! wl<355>   mc
XI833 blb vddh! wl<280>   mc
XI562 br vddh! wl<177>   mc
XI660 blb vddh! wl<488>   mc
XI570 brb vddh! wl<146>   mc
XI538 br vddh! wl<173>   mc
XI548 brb vddh! wl<184>   mc
XI529 brb vddh! wl<232>   mc
XI708 bl vddh! wl<451>   mc
XI668 blb vddh! wl<480>   mc
XI733 bl vddh! wl<325>   mc
XI756 bl vddh! wl<371>   mc
XI549 br vddh! wl<185>   mc
XI805 bl vddh! wl<313>   mc
XI551 brb vddh! wl<190>   mc
XI779 bl vddh! wl<365>   mc
XI539 brb vddh! wl<162>   mc
XI550 brb vddh! wl<186>   mc
XI530 br vddh! wl<235>   mc
XI563 br vddh! wl<145>   mc
XI612 blb vddh! wl<408>   mc
XI571 br vddh! wl<157>   mc
XI724 blb vddh! wl<328>   mc
XI652 bl vddh! wl<431>   mc
XI717 blb vddh! wl<460>   mc
XI764 bl vddh! wl<383>   mc
XI545 br vddh! wl<163>   mc
XI787 bl vddh! wl<299>   mc
XI536 brb vddh! wl<172>   mc
XI544 brb vddh! wl<166>   mc
XI527 brb vddh! wl<234>   mc
XI684 blb vddh! wl<496>   mc
XI693 blb vddh! wl<470>   mc
XI561 br vddh! wl<179>   mc
XI644 bl vddh! wl<419>   mc
XI569 brb vddh! wl<144>   mc
XI537 br vddh! wl<175>   mc
XI546 br vddh! wl<161>   mc
XI528 br vddh! wl<233>   mc
XI740 blb vddh! wl<344>   mc
XI547 br vddh! wl<187>   mc
XI796 blb vddh! wl<288>   mc
XI560 brb vddh! wl<182>   mc
XI568 br vddh! wl<149>   mc
XI700 bl vddh! wl<479>   mc
XI827 bl vddh! wl<285>   mc
XI677 bl vddh! wl<505>   mc
XI566 brb vddh! wl<148>   mc
XI557 br vddh! wl<181>   mc
XI629 blb vddh! wl<438>   mc
XI542 br vddh! wl<167>   mc
XI716 bl vddh! wl<463>   mc
XI533 br vddh! wl<169>   mc
XI685 bl vddh! wl<501>   mc
XI556 brb vddh! wl<176>   mc
XI573 brb vddh! wl<156>   mc
XI816 blb vddh! wl<310>   mc
XI732 blb vddh! wl<320>   mc
XI798 bl vddh! wl<295>   mc
XI849 blb vddh! wl<264>   mc
XI676 blb vddh! wl<504>   mc
XI543 brb vddh! wl<164>   mc
XI692 bl vddh! wl<467>   mc
XI534 brb vddh! wl<170>   mc
XI701 blb vddh! wl<476>   mc
XI558 br vddh! wl<183>   mc
XI574 brb vddh! wl<158>   mc
XI553 br vddh! wl<191>   mc
XI781 blb vddh! wl<364>   mc
XI540 brb vddh! wl<160>   mc
XI552 brb vddh! wl<188>   mc
XI531 br vddh! wl<171>   mc
XI709 blb vddh! wl<454>   mc
XI554 br vddh! wl<189>   mc
XI605 bl vddh! wl<389>   mc
XI565 brb vddh! wl<150>   mc
XI555 brb vddh! wl<178>   mc
XI541 br vddh! wl<165>   mc
XI532 brb vddh! wl<168>   mc
XI837 blb vddh! wl<262>   mc
XI620 blb vddh! wl<400>   mc
XI807 blb vddh! wl<318>   mc
XI564 br vddh! wl<147>   mc
XI604 blb vddh! wl<384>   mc
XI572 br vddh! wl<159>   mc
XI725 bl vddh! wl<329>   mc
XI628 bl vddh! wl<435>   mc
XI621 bl vddh! wl<405>   mc
XI690 bl vddh! wl<497>   mc
XI754 bl vddh! wl<337>   mc
XI516 br vddh! wl<227>   mc
XI730 bl vddh! wl<333>   mc
XI524 br vddh! wl<239>   mc
XI691 bl vddh! wl<465>   mc
XI507 br vddh! wl<253>   mc
XI486 brb vddh! wl<218>   mc
XI493 br vddh! wl<213>   mc
XI506 brb vddh! wl<242>   mc
XI659 bl vddh! wl<491>   mc
XI517 brb vddh! wl<230>   mc
XI618 bl vddh! wl<413>   mc
XI525 brb vddh! wl<236>   mc
XI714 blb vddh! wl<450>   mc
XI738 bl vddh! wl<321>   mc
XI492 brb vddh! wl<208>   mc
XI504 br vddh! wl<245>   mc
XI667 blb vddh! wl<482>   mc
XI731 blb vddh! wl<322>   mc
XI505 brb vddh! wl<240>   mc
XI485 br vddh! wl<217>   mc
XI847 blb vddh! wl<266>   mc
XI510 brb vddh! wl<254>   mc
XI746 bl vddh! wl<349>   mc
XI495 brb vddh! wl<212>   mc
XI626 bl vddh! wl<401>   mc
XI611 bl vddh! wl<411>   mc
XI699 bl vddh! wl<477>   mc
XI610 bl vddh! wl<385>   mc
XI675 bl vddh! wl<507>   mc
XI487 brb vddh! wl<222>   mc
XI825 blb vddh! wl<272>   mc
XI602 bl vddh! wl<397>   mc
XI762 blb vddh! wl<370>   mc
XI494 br vddh! wl<215>   mc
XI508 br vddh! wl<255>   mc
XI651 bl vddh! wl<429>   mc
XI518 brb vddh! wl<228>   mc
XI509 brb vddh! wl<252>   mc
XI526 brb vddh! wl<238>   mc
XI650 blb vddh! wl<418>   mc
XI683 blb vddh! wl<498>   mc
XI814 bl vddh! wl<311>   mc
XI512 br vddh! wl<249>   mc
XI707 bl vddh! wl<449>   mc
XI520 br vddh! wl<229>   mc
XI499 br vddh! wl<241>   mc
XI482 br vddh! wl<193>   mc
XI603 blb vddh! wl<386>   mc
XI498 br vddh! wl<209>   mc
XI513 brb vddh! wl<248>   mc
XI722 bl vddh! wl<459>   mc
XI521 brb vddh! wl<224>   mc
XI658 bl vddh! wl<427>   mc
XI723 bl vddh! wl<331>   mc
XI835 bl vddh! wl<257>   mc
XI627 bl vddh! wl<433>   mc
XI496 brb vddh! wl<214>   mc
XI826 blb vddh! wl<274>   mc
XI489 br vddh! wl<223>   mc
XI497 br vddh! wl<211>   mc
XI481 br vddh! wl<195>   mc
XI642 bl vddh! wl<443>   mc
XI698 blb vddh! wl<466>   mc
XI515 br vddh! wl<225>   mc
XI674 bl vddh! wl<481>   mc
XI523 br vddh! wl<237>   mc
XI491 brb vddh! wl<210>   mc
XI502 brb vddh! wl<244>   mc
XI643 bl vddh! wl<417>   mc
XI715 bl vddh! wl<461>   mc
XI503 br vddh! wl<247>   mc
XI484 brb vddh! wl<216>   mc
XI619 blb vddh! wl<402>   mc
XI501 brb vddh! wl<246>   mc
XI483 br vddh! wl<219>   mc
XI666 bl vddh! wl<493>   mc
XI706 bl vddh! wl<475>   mc
XI490 br vddh! wl<221>   mc
XI500 br vddh! wl<243>   mc
XI514 br vddh! wl<251>   mc
XI682 bl vddh! wl<509>   mc
XI522 brb vddh! wl<226>   mc
XI713 blb vddh! wl<448>   mc
XI770 bl vddh! wl<379>   mc
XI702 blb vddh! wl<478>   mc
XI729 bl vddh! wl<335>   mc
XI744 blb vddh! wl<348>   mc
XI649 blb vddh! wl<416>   mc
XI829 blb vddh! wl<284>   mc
XI760 bl vddh! wl<373>   mc
XI678 blb vddh! wl<506>   mc
XI818 bl vddh! wl<305>   mc
XI820 bl vddh! wl<275>   mc
XI734 bl vddh! wl<327>   mc
XI694 blb vddh! wl<468>   mc
XI705 blb vddh! wl<472>   mc
XI832 bl vddh! wl<281>   mc
XI689 bl vddh! wl<499>   mc
XI841 blb vddh! wl<256>   mc
XI670 bl vddh! wl<487>   mc
XI783 blb vddh! wl<362>   mc
XI726 blb vddh! wl<330>   mc
XI840 bl vddh! wl<261>   mc
XI822 blb vddh! wl<276>   mc
XI615 blb vddh! wl<414>   mc
XI679 blb vddh! wl<510>   mc
XI669 bl vddh! wl<485>   mc
XI804 blb vddh! wl<312>   mc
XI632 bl vddh! wl<437>   mc
XI703 blb vddh! wl<474>   mc
XI322 br vddh! wl<1>   mc
XI371 br vddh! wl<49>   mc
XI819 bl vddh! wl<273>   mc
XI321 br vddh! wl<3>   mc
XI782 blb vddh! wl<366>   mc
XI594 br vddh! wl<139>   mc
XI808 blb vddh! wl<316>   mc
XI593 brb vddh! wl<136>   mc
XI799 blb vddh! wl<292>   mc
XI592 br vddh! wl<137>   mc
XI790 blb vddh! wl<298>   mc
XI591 brb vddh! wl<138>   mc
XI749 bl vddh! wl<341>   mc
XI590 brb vddh! wl<142>   mc
XI765 blb vddh! wl<380>   mc
XI403 br vddh! wl<107>   mc
XI405 br vddh! wl<105>   mc
XI406 brb vddh! wl<106>   mc
XI407 brb vddh! wl<110>   mc
XI408 brb vddh! wl<108>   mc
XI409 br vddh! wl<111>   mc
XI411 brb vddh! wl<98>   mc
XI410 br vddh! wl<109>   mc
XI412 brb vddh! wl<96>   mc
XI413 br vddh! wl<101>   mc
XI414 br vddh! wl<103>   mc
XI415 brb vddh! wl<100>   mc
XI416 brb vddh! wl<102>   mc
XI417 br vddh! wl<99>   mc
XI418 br vddh! wl<97>   mc
XI420 brb vddh! wl<120>   mc
XI419 br vddh! wl<123>   mc
XI422 brb vddh! wl<122>   mc
XI421 br vddh! wl<121>   mc
XI423 brb vddh! wl<126>   mc
XI424 brb vddh! wl<124>   mc
XI425 br vddh! wl<127>   mc
XI426 br vddh! wl<125>   mc
XI427 brb vddh! wl<114>   mc
XI428 brb vddh! wl<112>   mc
XI429 br vddh! wl<117>   mc
XI430 br vddh! wl<119>   mc
XI402 br vddh! wl<43>   mc
XI401 brb vddh! wl<40>   mc
XI400 br vddh! wl<41>   mc
XI399 brb vddh! wl<42>   mc
XI398 brb vddh! wl<46>   mc
XI397 brb vddh! wl<44>   mc
XI310 brb vddh! wl<10>   mc
XI431 brb vddh! wl<116>   mc
XI396 br vddh! wl<47>   mc
XI801 bl vddh! wl<291>   mc
XI784 bl vddh! wl<361>   mc
XI395 br vddh! wl<45>   mc
XI735 blb vddh! wl<324>   mc
XI768 bl vddh! wl<377>   mc
XI663 blb vddh! wl<494>   mc
XI695 bl vddh! wl<471>   mc
XI759 bl vddh! wl<375>   mc
XI317 br vddh! wl<5>   mc
XI319 brb vddh! wl<4>   mc
XI600 blb vddh! wl<396>   mc
XI601 bl vddh! wl<399>   mc
XI655 blb vddh! wl<426>   mc
XI846 blb vddh! wl<270>   mc
XI751 blb vddh! wl<340>   mc
XI834 bl vddh! wl<283>   mc
XI743 blb vddh! wl<350>   mc
XI719 blb vddh! wl<458>   mc
XI792 blb vddh! wl<300>   mc
XI671 blb vddh! wl<484>   mc
XI623 blb vddh! wl<404>   mc
XI810 bl vddh! wl<317>   mc
XI647 bl vddh! wl<423>   mc
XI780 bl vddh! wl<367>   mc
XI475 brb vddh! wl<194>   mc
XI635 bl vddh! wl<445>   mc
XI467 br vddh! wl<203>   mc
XI771 bl vddh! wl<353>   mc
XI769 blb vddh! wl<376>   mc
XI806 blb vddh! wl<314>   mc
XI476 brb vddh! wl<192>   mc
XI633 blb vddh! wl<432>   mc
XI394 brb vddh! wl<34>   mc
XI393 brb vddh! wl<32>   mc
XI468 brb vddh! wl<200>   mc
XI803 bl vddh! wl<315>   mc
XI794 bl vddh! wl<301>   mc
XI392 br vddh! wl<37>   mc
XI391 br vddh! wl<39>   mc
XI474 br vddh! wl<205>   mc
XI390 brb vddh! wl<36>   mc
XI774 blb vddh! wl<356>   mc
XI755 bl vddh! wl<369>   mc
XI307 br vddh! wl<11>   mc
XI824 bl vddh! wl<277>   mc
XI389 brb vddh! wl<38>   mc
XI795 blb vddh! wl<290>   mc
XI812 blb vddh! wl<304>   mc
XI388 br vddh! wl<35>   mc
XI320 brb vddh! wl<6>   mc
XI387 br vddh! wl<33>   mc
XI598 blb vddh! wl<394>   mc
XI386 br vddh! wl<59>   mc
XI385 brb vddh! wl<56>   mc
XI384 br vddh! wl<57>   mc
XI383 brb vddh! wl<58>   mc
XI381 brb vddh! wl<60>   mc
XI382 brb vddh! wl<62>   mc
XI380 br vddh! wl<63>   mc
XI379 br vddh! wl<61>   mc
XI378 brb vddh! wl<50>   mc
XI377 brb vddh! wl<48>   mc
XI599 blb vddh! wl<398>   mc
XI376 br vddh! wl<53>   mc
XI375 br vddh! wl<55>   mc
XI773 blb vddh! wl<358>   mc
XI374 brb vddh! wl<52>   mc
XI373 brb vddh! wl<54>   mc
XI372 br vddh! wl<51>   mc
XI711 bl vddh! wl<455>   mc
XI786 bl vddh! wl<363>   mc
XI687 blb vddh! wl<500>   mc
XI830 blb vddh! wl<286>   mc
XI739 bl vddh! wl<347>   mc
XI637 blb vddh! wl<444>   mc
XI432 brb vddh! wl<118>   mc
XI638 blb vddh! wl<446>   mc
XI473 br vddh! wl<207>   mc
XI433 br vddh! wl<115>   mc
XI775 bl vddh! wl<359>   mc
XI848 bl vddh! wl<265>   mc
XI641 blb vddh! wl<440>   mc
XI747 blb vddh! wl<338>   mc
XI479 brb vddh! wl<196>   mc
XI823 bl vddh! wl<279>   mc
XI471 brb vddh! wl<206>   mc
XI778 blb vddh! wl<354>   mc
XI844 bl vddh! wl<271>   mc
XI776 bl vddh! wl<357>   mc
XI313 br vddh! wl<15>   mc
XI777 blb vddh! wl<352>   mc
XI434 br vddh! wl<113>   mc
XI435 br vddh! wl<81>   mc
XI480 brb vddh! wl<198>   mc
XI640 bl vddh! wl<441>   mc
XI472 brb vddh! wl<204>   mc
XI767 blb vddh! wl<378>   mc
XI478 br vddh! wl<199>   mc
XI311 brb vddh! wl<14>   mc
XI309 br vddh! wl<9>   mc
XI843 bl vddh! wl<269>   mc
XI314 br vddh! wl<13>   mc
XI470 brb vddh! wl<202>   mc
XI436 br vddh! wl<83>   mc
XI815 blb vddh! wl<308>   mc
XI323 br vddh! wl<27>   mc
XI437 brb vddh! wl<86>   mc
XI788 blb vddh! wl<296>   mc
XI438 brb vddh! wl<84>   mc
XI439 br vddh! wl<87>   mc
XI440 br vddh! wl<85>   mc
XI441 brb vddh! wl<80>   mc
XI442 brb vddh! wl<82>   mc
XI845 blb vddh! wl<268>   mc
XI836 bl vddh! wl<259>   mc
XI797 bl vddh! wl<293>   mc
XI443 br vddh! wl<93>   mc
XI477 br vddh! wl<197>   mc
XI631 bl vddh! wl<439>   mc
XI469 br vddh! wl<201>   mc
XI681 bl vddh! wl<511>   mc
XI821 blb vddh! wl<278>   mc
XI648 bl vddh! wl<421>   mc
XI697 blb vddh! wl<464>   mc
XI315 brb vddh! wl<2>   mc
XI606 bl vddh! wl<391>   mc
XI656 bl vddh! wl<425>   mc
XI758 blb vddh! wl<372>   mc
XI672 blb vddh! wl<486>   mc
XI444 br vddh! wl<95>   mc
XI445 brb vddh! wl<92>   mc
XI324 brb vddh! wl<24>   mc
XI325 br vddh! wl<25>   mc
XI326 brb vddh! wl<26>   mc
XI446 brb vddh! wl<94>   mc
XI447 brb vddh! wl<90>   mc
XI327 brb vddh! wl<30>   mc
XI448 br vddh! wl<89>   mc
XI328 brb vddh! wl<28>   mc
XI616 blb vddh! wl<412>   mc
XI329 br vddh! wl<31>   mc
XI449 brb vddh! wl<88>   mc
XI450 br vddh! wl<91>   mc
XI451 br vddh! wl<65>   mc
XI452 br vddh! wl<67>   mc
XI453 brb vddh! wl<70>   mc
XI454 brb vddh! wl<68>   mc
XI721 blb vddh! wl<456>   mc
XI842 blb vddh! wl<258>   mc
XI664 blb vddh! wl<492>   mc
XI737 bl vddh! wl<323>   mc
XI718 blb vddh! wl<462>   mc
XI831 blb vddh! wl<282>   mc
XI839 bl vddh! wl<263>   mc
XI622 bl vddh! wl<407>   mc
XI455 br vddh! wl<71>   mc
XI745 bl vddh! wl<351>   mc
XI736 blb vddh! wl<326>   mc
XI609 bl vddh! wl<387>   mc
XI330 br vddh! wl<29>   mc
XI331 brb vddh! wl<18>   mc
XI404 brb vddh! wl<104>   mc
XI316 brb vddh! wl<0>   mc
XI654 blb vddh! wl<430>   mc
XI720 bl vddh! wl<457>   mc
XI750 bl vddh! wl<343>   mc
XI696 bl vddh! wl<469>   mc
XI332 brb vddh! wl<16>   mc
XI791 blb vddh! wl<302>   mc
XI614 blb vddh! wl<410>   mc
XI595 bl vddh! wl<395>   mc
XI608 blb vddh! wl<390>   mc
XI333 br vddh! wl<21>   mc
XI308 brb vddh! wl<8>   mc
XI766 blb vddh! wl<382>   mc
XI456 br vddh! wl<69>   mc
XI625 bl vddh! wl<403>   mc
XI596 blb vddh! wl<392>   mc
XI597 bl vddh! wl<393>   mc
XI630 blb vddh! wl<436>   mc
XI634 blb vddh! wl<434>   mc
XI457 brb vddh! wl<64>   mc
XI742 blb vddh! wl<346>   mc
XI761 blb vddh! wl<368>   mc
XI318 br vddh! wl<7>   mc
XI624 blb vddh! wl<406>   mc
XI617 bl vddh! wl<415>   mc
XI809 bl vddh! wl<319>   mc
XI458 brb vddh! wl<66>   mc
XI459 br vddh! wl<77>   mc
XI460 br vddh! wl<79>   mc
XI334 br vddh! wl<23>   mc
XI704 bl vddh! wl<473>   mc
XI657 blb vddh! wl<424>   mc
XI785 blb vddh! wl<360>   mc
XI335 brb vddh! wl<20>   mc
XI461 brb vddh! wl<76>   mc
XI688 blb vddh! wl<502>   mc
XI336 brb vddh! wl<22>   mc
XI337 br vddh! wl<19>   mc
XI686 bl vddh! wl<503>   mc
XI793 bl vddh! wl<303>   mc
XI462 brb vddh! wl<78>   mc
XI338 br vddh! wl<17>   mc
XI710 blb vddh! wl<452>   mc
XI463 brb vddh! wl<74>   mc
XI811 blb vddh! wl<306>   mc
XI646 blb vddh! wl<420>   mc
XI673 bl vddh! wl<483>   mc
XI752 blb vddh! wl<342>   mc
XI728 blb vddh! wl<332>   mc
XI464 br vddh! wl<73>   mc
XI665 bl vddh! wl<495>   mc
XI802 bl vddh! wl<289>   mc
XI712 bl vddh! wl<453>   mc
XI312 brb vddh! wl<12>   mc
XI465 brb vddh! wl<72>   mc
XI466 br vddh! wl<75>   mc
XI727 blb vddh! wl<334>   mc
XI800 blb vddh! wl<294>   mc
XI304 bl blb br brb cs io io_ l_sel n_ena p_ena pre r_sel   sa_pre
CC51 blb gnd! 250f $[CP]
CC52 bl gnd! 250f $[CP]
CC8 brb gnd! 250f $[CP]
CC7 br gnd! 250f $[CP]
.ENDS
