.SUBCKT decoder4_16 A<3> A<2> A<1> A<0> ENA X<15> X<14> X<13> X<12> X<11>
+X<10> X<9> X<8> X<7> X<6> X<5> X<4> X<3> X<2> X<1> X<0>
XI27 net146 net142 net138 net132 net128 net126   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI17 net146 net117 net138 net134 net128 net131   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI32 net146 net142 net136 net132 net130 net286   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI31 net146 net142 net136 net132 net128 net285   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI30 net146 net142 net136 net134 net130 net150   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI29 net146 net142 net136 net134 net128 net156   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI23 net146 net117 net136 net132 net128 net162   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI19 net146 net117 net138 net132 net128 net168   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI24 net146 net117 net136 net132 net130 net174   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI20 net146 net117 net138 net132 net130 net180   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI21 net146 net117 net136 net134 net128 net186   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI22 net146 net117 net136 net134 net130 net192   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI18 net146 net117 net138 net134 net130 net198   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI26 net146 net142 net138 net134 net130 net204   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI28 net146 net142 net138 net132 net130 net210   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI25 net146 net142 net138 net134 net128 net216   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI93 ENA net144   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=4.2u
XI45 net198 X<14>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI46 net168 X<13>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI47 net180 X<12>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI44 net131 X<15>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI48 net186 X<11>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI49 net192 X<10>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI50 net162 X<9>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI51 net174 X<8>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI52 net216 X<7>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI53 net204 X<6>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI54 net126 X<5>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI55 net210 X<4>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI56 net156 X<3>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI57 net150 X<2>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI58 net285 X<1>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI59 net286 X<0>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI42 net144 net146   inv Ln=0.35u Wn=2.1u M=3 Lp=0.35u Wp=4.2u
XI41 A<1> net132   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=3.2u
XI40 net132 net134   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=3.2u
XI39 net130 net128   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=3.2u
XI38 A<0> net130   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=3.2u
XI37 A<2> net136   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=3.2u
XI33 A<3> net142   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=3.2u
XI36 net136 net138   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=3.2u
XI35 net142 net117   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=3.2u
.ENDS
