.SUBCKT atd18 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7>
+a<6> a<5> a<4> a<3> a<2> a<1> a<0> w_ y
XI103 net99 net97 net189 net163   nor3 Lp=0.35u Wp=7u Ln=0.35u Wn=3.5u
XI74 net157 net152 net147 net142 net163 net137   nand5 Lp=0.35u Wp=4u Ln=0.35u
+Wn=7u
XI96 net169 net165 net171 net167 net142   nor4 Lp=0.35u Wp=7u Ln=0.35u Wn=3.5u
XI93 net181 net183 net187 net185 net152   nor4 Lp=0.35u Wp=7u Ln=0.35u Wn=3.5u
XI92 net193 net195 net197 net191 net157   nor4 Lp=0.35u Wp=7u Ln=0.35u Wn=3.5u
XI94 net175 net179 net173 net177 net147   nor4 Lp=0.35u Wp=7u Ln=0.35u Wn=3.5u
XI75 net137 net159   inv Ln=0.35u Wn=8u M=3 Lp=0.35u Wp=16u
XI81 net159 y   inv Ln=0.35u Wn=8u M=9 Lp=0.35u Wp=16u
XI101 a<16> net99   atd1
XI102 a<17> net97   atd1
XI97 a<14> net171   atd1
XI98 a<12> net169   atd1
XI71 a<3> net191   atd1
XI99 a<15> net167   atd1
XI79 w_ net189   atd1
XI91 a<10> net173   atd1
XI68 a<0> net193   atd1
XI83 a<4> net181   atd1
XI84 a<5> net183   atd1
XI82 a<7> net185   atd1
XI88 a<8> net175   atd1
XI85 a<6> net187   atd1
XI100 a<13> net165   atd1
XI69 a<1> net195   atd1
XI70 a<2> net197   atd1
XI90 a<11> net177   atd1
XI89 a<9> net179   atd1
.ENDS
