.SUBCKT io a0 i_o io io_ main_ena pre w_
MM0 net52 net107 gnd! vbb! NMOS W=1.4u L=350.00n M=1
MM12 i_o net93 net52 vbb! NMOS W=1.4u L=350.00n M=1
MM1 i_o net101 net63 vdd! PMOS W=3.5u L=350.00n M=1
MM2 net63 net107 vdd! vdd! PMOS W=3.5u L=350.00n M=1
XI210 main_ena io io_ net73 net70 pre   main_sense
XI218 net73 net83 net111 a0   ctg Lp=0.35u Wp=3.5u Ln=0.35u Wn=3.5u
XI196 io_ net95 a0 net119   ctg Lp=0.35u Wp=3.5u Ln=0.35u Wn=3.5u
XI164 io net95 net119 a0   ctg Lp=0.35u Wp=3.5u Ln=0.35u Wn=3.5u
XI161 net95 i_o net101 net93   ctg Lp=0.35u Wp=3.5u Ln=0.35u Wn=3.5u
XI217 net70 net83 a0 net111   ctg Lp=0.35u Wp=3.5u Ln=0.35u Wn=3.5u
XI224 net83 net107   inv Ln=0.35u Wn=1.4u M=1 Lp=0.35u Wp=2.8u
XI306 w_ net101   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI165 a0 net119   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI307 net101 net93   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI219 a0 net111   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI195 io io_ pre   precharge
CC20 io_ gnd! 200f $[CP]
CC22 io gnd! 200f $[CP]
.ENDS
