.SUBCKT block512x512n a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9>
+a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> ena i_o w_
XI102 net696 i_o ena net690   ctg Lp=0.35u Wp=1.4u Ln=0.35u Wn=1.4u
XI100 ena net690   inv Ln=0.35u Wn=1.4u M=1 Lp=0.35u Wp=1.4u
XI1367 a<0> net696 net9403 net9404 main_ena pre w_   io
XI1366 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6>
+a<5> a<4> a<3> a<2> a<1> a<0> cl<511> cl<510> cl<509> cl<508> cl<507> cl<506>
+cl<505> cl<504> cl<503> cl<502> cl<501> cl<500> cl<499> cl<498> cl<497>
+cl<496> cl<495> cl<494> cl<493> cl<492> cl<491> cl<490> cl<489> cl<488>
+cl<487> cl<486> cl<485> cl<484> cl<483> cl<482> cl<481> cl<480> cl<479>
+cl<478> cl<477> cl<476> cl<475> cl<474> cl<473> cl<472> cl<471> cl<470>
+cl<469> cl<468> cl<467> cl<466> cl<465> cl<464> cl<463> cl<462> cl<461>
+cl<460> cl<459> cl<458> cl<457> cl<456> cl<455> cl<454> cl<453> cl<452>
+cl<451> cl<450> cl<449> cl<448> cl<447> cl<446> cl<445> cl<444> cl<443>
+cl<442> cl<441> cl<440> cl<439> cl<438> cl<437> cl<436> cl<435> cl<434>
+cl<433> cl<432> cl<431> cl<430> cl<429> cl<428> cl<427> cl<426> cl<425>
+cl<424> cl<423> cl<422> cl<421> cl<420> cl<419> cl<418> cl<417> cl<416>
+cl<415> cl<414> cl<413> cl<412> cl<411> cl<410> cl<409> cl<408> cl<407>
+cl<406> cl<405> cl<404> cl<403> cl<402> cl<401> cl<400> cl<399> cl<398>
+cl<397> cl<396> cl<395> cl<394> cl<393> cl<392> cl<391> cl<390> cl<389>
+cl<388> cl<387> cl<386> cl<385> cl<384> cl<383> cl<382> cl<381> cl<380>
+cl<379> cl<378> cl<377> cl<376> cl<375> cl<374> cl<373> cl<372> cl<371>
+cl<370> cl<369> cl<368> cl<367> cl<366> cl<365> cl<364> cl<363> cl<362>
+cl<361> cl<360> cl<359> cl<358> cl<357> cl<356> cl<355> cl<354> cl<353>
+cl<352> cl<351> cl<350> cl<349> cl<348> cl<347> cl<346> cl<345> cl<344>
+cl<343> cl<342> cl<341> cl<340> cl<339> cl<338> cl<337> cl<336> cl<335>
+cl<334> cl<333> cl<332> cl<331> cl<330> cl<329> cl<328> cl<327> cl<326>
+cl<325> cl<324> cl<323> cl<322> cl<321> cl<320> cl<319> cl<318> cl<317>
+cl<316> cl<315> cl<314> cl<313> cl<312> cl<311> cl<310> cl<309> cl<308>
+cl<307> cl<306> cl<305> cl<304> cl<303> cl<302> cl<301> cl<300> cl<299>
+cl<298> cl<297> cl<296> cl<295> cl<294> cl<293> cl<292> cl<291> cl<290>
+cl<289> cl<288> cl<287> cl<286> cl<285> cl<284> cl<283> cl<282> cl<281>
+cl<280> cl<279> cl<278> cl<277> cl<276> cl<275> cl<274> cl<273> cl<272>
+cl<271> cl<270> cl<269> cl<268> cl<267> cl<266> cl<265> cl<264> cl<263>
+cl<262> cl<261> cl<260> cl<259> cl<258> cl<257> cl<256> cl<255> cl<254>
+cl<253> cl<252> cl<251> cl<250> cl<249> cl<248> cl<247> cl<246> cl<245>
+cl<244> cl<243> cl<242> cl<241> cl<240> cl<239> cl<238> cl<237> cl<236>
+cl<235> cl<234> cl<233> cl<232> cl<231> cl<230> cl<229> cl<228> cl<227>
+cl<226> cl<225> cl<224> cl<223> cl<222> cl<221> cl<220> cl<219> cl<218>
+cl<217> cl<216> cl<215> cl<214> cl<213> cl<212> cl<211> cl<210> cl<209>
+cl<208> cl<207> cl<206> cl<205> cl<204> cl<203> cl<202> cl<201> cl<200>
+cl<199> cl<198> cl<197> cl<196> cl<195> cl<194> cl<193> cl<192> cl<191>
+cl<190> cl<189> cl<188> cl<187> cl<186> cl<185> cl<184> cl<183> cl<182>
+cl<181> cl<180> cl<179> cl<178> cl<177> cl<176> cl<175> cl<174> cl<173>
+cl<172> cl<171> cl<170> cl<169> cl<168> cl<167> cl<166> cl<165> cl<164>
+cl<163> cl<162> cl<161> cl<160> cl<159> cl<158> cl<157> cl<156> cl<155>
+cl<154> cl<153> cl<152> cl<151> cl<150> cl<149> cl<148> cl<147> cl<146>
+cl<145> cl<144> cl<143> cl<142> cl<141> cl<140> cl<139> cl<138> cl<137>
+cl<136> cl<135> cl<134> cl<133> cl<132> cl<131> cl<130> cl<129> cl<128>
+cl<127> cl<126> cl<125> cl<124> cl<123> cl<122> cl<121> cl<120> cl<119>
+cl<118> cl<117> cl<116> cl<115> cl<114> cl<113> cl<112> cl<111> cl<110>
+cl<109> cl<108> cl<107> cl<106> cl<105> cl<104> cl<103> cl<102> cl<101>
+cl<100> cl<99> cl<98> cl<97> cl<96> cl<95> cl<94> cl<93> cl<92> cl<91> cl<90>
+cl<89> cl<88> cl<87> cl<86> cl<85> cl<84> cl<83> cl<82> cl<81> cl<80> cl<79>
+cl<78> cl<77> cl<76> cl<75> cl<74> cl<73> cl<72> cl<71> cl<70> cl<69> cl<68>
+cl<67> cl<66> cl<65> cl<64> cl<63> cl<62> cl<61> cl<60> cl<59> cl<58> cl<57>
+cl<56> cl<55> cl<54> cl<53> cl<52> cl<51> cl<50> cl<49> cl<48> cl<47> cl<46>
+cl<45> cl<44> cl<43> cl<42> cl<41> cl<40> cl<39> cl<38> cl<37> cl<36> cl<35>
+cl<34> cl<33> cl<32> cl<31> cl<30> cl<29> cl<28> cl<27> cl<26> cl<25> cl<24>
+cl<23> cl<22> cl<21> cl<20> cl<19> cl<18> cl<17> cl<16> cl<15> cl<14> cl<13>
+cl<12> cl<11> cl<10> cl<9> cl<8> cl<7> cl<6> cl<5> cl<4> cl<3> cl<2> cl<1>
+cl<0> ena l_sel main_ena n_ena p_ena pre r_sel w_ wl<511> wl<510> wl<509>
+wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501> wl<500>
+wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492> wl<491>
+wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483> wl<482>
+wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474> wl<473>
+wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465> wl<464>
+wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456> wl<455>
+wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447> wl<446>
+wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438> wl<437>
+wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429> wl<428>
+wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420> wl<419>
+wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411> wl<410>
+wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402> wl<401>
+wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393> wl<392>
+wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384> wl<383>
+wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375> wl<374>
+wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366> wl<365>
+wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357> wl<356>
+wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348> wl<347>
+wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339> wl<338>
+wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330> wl<329>
+wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321> wl<320>
+wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312> wl<311>
+wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303> wl<302>
+wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294> wl<293>
+wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285> wl<284>
+wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276> wl<275>
+wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267> wl<266>
+wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258> wl<257>
+wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249> wl<248>
+wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240> wl<239>
+wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231> wl<230>
+wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222> wl<221>
+wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213> wl<212>
+wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204> wl<203>
+wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195> wl<194>
+wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186> wl<185>
+wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177> wl<176>
+wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168> wl<167>
+wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159> wl<158>
+wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150> wl<149>
+wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141> wl<140>
+wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132> wl<131>
+wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123> wl<122>
+wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114> wl<113>
+wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105> wl<104>
+wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95> wl<94>
+wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84> wl<83>
+wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73> wl<72>
+wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62> wl<61>
+wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51> wl<50>
+wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40> wl<39>
+wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29> wl<28>
+wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18> wl<17>
+wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7> wl<6>
+wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   ctrl256kbm
XI887 cl<34> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI888 cl<38> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI889 cl<44> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI890 cl<39> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI891 cl<37> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI892 cl<36> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI893 cl<45> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI894 cl<47> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI895 cl<46> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI896 cl<42> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI897 cl<43> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI898 cl<41> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI899 cl<40> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI900 cl<56> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI901 cl<57> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI902 cl<59> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI903 cl<58> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI904 cl<62> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI905 cl<63> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI906 cl<61> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI907 cl<60> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI908 cl<52> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI909 cl<53> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI910 cl<55> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI911 cl<54> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI912 cl<50> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI913 cl<51> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI914 cl<49> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI915 cl<48> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI916 cl<32> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI917 cl<33> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI918 cl<97> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI919 cl<96> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI920 cl<112> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI922 cl<115> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI923 cl<114> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI921 cl<113> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI924 cl<118> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI925 cl<119> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI926 cl<117> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI927 cl<116> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI928 cl<124> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI929 cl<125> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI930 cl<127> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI931 cl<126> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI932 cl<122> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI933 cl<123> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI934 cl<121> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI935 cl<120> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI936 cl<104> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI937 cl<105> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI938 cl<107> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI939 cl<106> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI940 cl<110> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI941 cl<111> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI942 cl<109> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI943 cl<100> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI944 cl<101> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI945 cl<103> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI946 cl<108> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI947 cl<102> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI948 cl<98> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI949 cl<99> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI950 cl<67> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI951 cl<66> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI952 cl<70> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI953 cl<76> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI954 cl<71> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI955 cl<69> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI956 cl<68> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI957 cl<77> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI958 cl<79> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI959 cl<78> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI960 cl<74> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI961 cl<75> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI962 cl<73> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI963 cl<72> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI964 cl<88> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI965 cl<89> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI966 cl<91> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI967 cl<90> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI968 cl<94> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI969 cl<95> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI970 cl<93> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI971 cl<92> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI972 cl<84> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI973 cl<85> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI974 cl<87> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI975 cl<86> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI976 cl<82> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI977 cl<83> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI978 cl<81> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI979 cl<80> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI980 cl<64> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI981 cl<65> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI982 cl<193> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI983 cl<192> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI984 cl<208> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI987 cl<210> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI988 cl<214> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI985 cl<209> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI986 cl<211> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI989 cl<215> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI990 cl<213> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI991 cl<212> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI992 cl<220> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI993 cl<221> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI994 cl<223> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI995 cl<222> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI996 cl<219> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI997 cl<218> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI998 cl<217> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI999 cl<216> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1000 cl<200> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1001 cl<201> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1002 cl<203> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1003 cl<202> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1004 cl<206> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1005 cl<207> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1006 cl<205> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1007 cl<196> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1008 cl<197> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1009 cl<199> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1010 cl<204> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1011 cl<198> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1012 cl<194> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1013 cl<195> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1014 cl<227> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1015 cl<226> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1016 cl<230> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1017 cl<236> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1018 cl<231> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1019 cl<229> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1020 cl<228> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1021 cl<237> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1022 cl<239> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1023 cl<238> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1024 cl<234> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1025 cl<235> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1026 cl<233> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1027 cl<232> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1028 cl<248> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1029 cl<249> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1030 cl<251> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1031 cl<250> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1032 cl<254> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1033 cl<255> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1034 cl<253> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1035 cl<252> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1036 cl<244> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1037 cl<245> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1038 cl<247> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1039 cl<246> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1040 cl<242> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1041 cl<243> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1042 cl<241> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1043 cl<240> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1044 cl<224> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1045 cl<225> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1046 cl<161> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1047 cl<160> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1048 cl<176> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1049 cl<177> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1050 cl<179> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1051 cl<178> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1052 cl<182> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1053 cl<183> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1054 cl<181> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1055 cl<180> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1056 cl<188> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1057 cl<189> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1058 cl<191> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1059 cl<190> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1060 cl<186> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1061 cl<187> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1062 cl<185> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1063 cl<184> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1064 cl<168> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1065 cl<169> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1066 cl<171> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1067 cl<170> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1068 cl<174> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1069 cl<175> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1070 cl<173> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1071 cl<164> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1072 cl<165> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1073 cl<167> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1074 cl<172> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1075 cl<166> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1076 cl<162> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1077 cl<163> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1078 cl<131> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1079 cl<130> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1080 cl<134> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1081 cl<140> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1082 cl<135> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1083 cl<133> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1084 cl<132> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1085 cl<141> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1086 cl<143> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1087 cl<142> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1088 cl<138> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1089 cl<139> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1090 cl<137> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1091 cl<136> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1092 cl<152> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1093 cl<153> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1094 cl<155> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1095 cl<154> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1096 cl<158> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1097 cl<159> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1098 cl<157> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1099 cl<156> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1100 cl<148> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1101 cl<149> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1102 cl<151> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1103 cl<150> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1104 cl<146> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1105 cl<147> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1106 cl<145> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1107 cl<144> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1108 cl<128> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1109 cl<129> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1110 cl<385> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1111 cl<384> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1114 cl<403> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI856 cl<3> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI857 cl<2> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI858 cl<6> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI862 cl<12> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI859 cl<7> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI860 cl<5> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI861 cl<4> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI863 cl<13> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI864 cl<15> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI865 cl<14> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI866 cl<10> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI867 cl<11> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI868 cl<9> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI869 cl<8> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI870 cl<24> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI871 cl<25> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI872 cl<27> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI873 cl<26> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI874 cl<30> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI875 cl<31> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI876 cl<29> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI877 cl<28> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI878 cl<20> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI879 cl<21> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI880 cl<23> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI881 cl<22> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI882 cl<18> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI883 cl<19> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI884 cl<17> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI885 cl<16> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1115 cl<402> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1112 cl<400> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1113 cl<401> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1116 cl<406> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1117 cl<407> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1118 cl<405> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1119 cl<404> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1120 cl<412> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1121 cl<413> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1122 cl<415> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1123 cl<414> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1124 cl<410> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1125 cl<411> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1126 cl<409> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1127 cl<408> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1128 cl<392> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1129 cl<393> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1130 cl<395> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1131 cl<394> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1132 cl<398> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1133 cl<399> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1134 cl<397> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1135 cl<388> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1136 cl<389> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1137 cl<391> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1138 cl<396> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1139 cl<390> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1140 cl<386> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1141 cl<387> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1142 cl<419> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1143 cl<418> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1144 cl<422> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1145 cl<428> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1146 cl<423> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1147 cl<421> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1148 cl<420> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1149 cl<429> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1150 cl<431> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1151 cl<430> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1152 cl<426> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1153 cl<427> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1154 cl<425> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1155 cl<424> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1156 cl<440> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1157 cl<441> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1158 cl<443> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1159 cl<442> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1160 cl<446> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1161 cl<447> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1162 cl<445> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1163 cl<444> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1164 cl<436> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1165 cl<437> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1166 cl<439> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1167 cl<438> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1168 cl<434> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1169 cl<435> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1170 cl<433> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1171 cl<432> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1172 cl<416> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1173 cl<417> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1174 cl<481> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1175 cl<480> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1176 cl<496> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1177 cl<497> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1178 cl<499> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1179 cl<498> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1180 cl<502> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1181 cl<503> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1182 cl<501> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1183 cl<500> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1184 cl<508> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1185 cl<509> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1186 cl<511> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1187 cl<510> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1188 cl<506> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1189 cl<507> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1190 cl<505> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1191 cl<504> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1192 cl<488> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1193 cl<489> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1194 cl<491> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1195 cl<490> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1196 cl<494> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1197 cl<495> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1198 cl<493> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1199 cl<484> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1200 cl<485> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1201 cl<487> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1202 cl<492> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1203 cl<486> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1204 cl<482> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1205 cl<483> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1206 cl<451> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1207 cl<450> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1208 cl<454> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1209 cl<460> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1210 cl<455> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1211 cl<453> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1212 cl<452> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1213 cl<461> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1214 cl<463> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1215 cl<462> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1216 cl<458> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1217 cl<459> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1218 cl<457> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1219 cl<456> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1220 cl<472> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1221 cl<473> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1222 cl<475> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1223 cl<474> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1224 cl<478> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1225 cl<479> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1226 cl<477> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1227 cl<476> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1228 cl<468> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1229 cl<469> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1230 cl<471> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1231 cl<470> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1232 cl<466> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1233 cl<467> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1234 cl<465> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1235 cl<464> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1236 cl<448> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1237 cl<449> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1238 cl<321> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1239 cl<320> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1240 cl<336> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1241 cl<337> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1242 cl<339> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1243 cl<338> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1244 cl<342> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1245 cl<343> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1246 cl<341> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1247 cl<340> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1248 cl<348> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1249 cl<349> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1250 cl<351> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1251 cl<350> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1252 cl<346> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1253 cl<347> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1254 cl<345> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1255 cl<344> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1256 cl<328> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1257 cl<329> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1258 cl<331> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1259 cl<330> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1260 cl<334> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1261 cl<335> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1262 cl<333> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1263 cl<324> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1264 cl<325> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1265 cl<327> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1266 cl<332> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1267 cl<326> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1268 cl<322> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1269 cl<323> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1270 cl<355> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1271 cl<354> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1272 cl<358> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1273 cl<364> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1274 cl<359> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1275 cl<357> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1276 cl<356> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1277 cl<365> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1278 cl<367> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1279 cl<366> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1280 cl<362> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1281 cl<363> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1282 cl<361> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1283 cl<360> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1284 cl<376> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1285 cl<377> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1286 cl<379> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1287 cl<378> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1288 cl<382> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1289 cl<383> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1290 cl<381> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1291 cl<380> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1292 cl<372> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1293 cl<373> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1294 cl<375> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1295 cl<374> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1296 cl<370> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1297 cl<371> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1298 cl<369> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1299 cl<368> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1300 cl<352> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1301 cl<353> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1302 cl<289> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1303 cl<288> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1304 cl<304> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1305 cl<305> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1306 cl<307> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1307 cl<306> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1308 cl<310> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1309 cl<311> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1310 cl<309> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1311 cl<308> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1312 cl<316> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1313 cl<317> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1314 cl<319> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1315 cl<318> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1316 cl<314> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1317 cl<315> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1318 cl<313> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1319 cl<312> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1320 cl<296> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1321 cl<297> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1322 cl<299> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1323 cl<298> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1324 cl<302> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1325 cl<303> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1326 cl<301> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1327 cl<292> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1328 cl<293> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1329 cl<295> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1330 cl<300> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1331 cl<294> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1332 cl<290> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1333 cl<291> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1334 cl<259> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1335 cl<258> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1336 cl<262> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1337 cl<268> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1338 cl<263> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1339 cl<261> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1340 cl<260> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1341 cl<269> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1342 cl<271> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1343 cl<270> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1344 cl<266> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1345 cl<267> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1346 cl<265> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1347 cl<264> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1348 cl<280> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1349 cl<281> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1350 cl<283> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1351 cl<282> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1352 cl<286> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1353 cl<287> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1354 cl<285> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1355 cl<284> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1356 cl<276> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1357 cl<277> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1358 cl<279> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1359 cl<278> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1360 cl<274> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1361 cl<275> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1362 cl<273> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1363 cl<272> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1364 cl<256> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1365 cl<257> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI886 cl<35> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI854 cl<0> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI855 cl<1> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
.ENDS
