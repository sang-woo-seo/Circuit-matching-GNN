.SUBCKT dram1gbn a<29> a<28> a<27> a<26> a<25> a<24> a<23> a<22> a<21> a<20>
+a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7>
+a<6> a<5> a<4> a<3> a<2> a<1> a<0> d ena q w_
XI66 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<22> 0 net230
+  bank16mx1n
XI65 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<6> 0 net230
+  bank16mx1n
XI64 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<23> 0 net230
+  bank16mx1n
XI63 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<7> 0 net230
+  bank16mx1n
XI62 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<8> 0 net230
+  bank16mx1n
XI61 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<25> 0 net230
+  bank16mx1n
XI59 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<27> 0 net230
+  bank16mx1n
XI58 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<24> 0 net230
+  bank16mx1n
***XI57 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<20> 0 net230
***+  bank16mx1n
***XI56 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<21> 0 net230
***+  bank16mx1n
***XI55 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<26> 0 net230
***+  bank16mx1n
***XI54 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<4> 0 net230
***+  bank16mx1n
***XI53 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<11> 0 net230
***+  bank16mx1n
***XI52 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<5> 0 net230
***+  bank16mx1n
***XI49 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<10> 0 net230
***+  bank16mx1n
***XI35 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<39> 0 net230
***+  bank16mx1n
***XI36 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<40> 0 net230
***+  bank16mx1n
***XI41 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<52> 0 net230
***+  bank16mx1n
***XI32 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<54> 0 net230
***+  bank16mx1n
***XI47 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<41> 0 net230
***+  bank16mx1n
***XI51 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<9> 0 net230
***+  bank16mx1n
***XI38 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<59> 0 net230
***+  bank16mx1n
***XI48 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<42> 0 net230
***+  bank16mx1n
***XI18 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<33> 0 net230
***+  bank16mx1n
***XI21 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<62> 0 net230
***+  bank16mx1n
***XI20 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<32> 0 net230
***+  bank16mx1n
***XI42 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<53> 0 net230
***+  bank16mx1n
***XI22 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<49> 0 net230
***+  bank16mx1n
***XI28 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<35> 0 net230
***+  bank16mx1n
***XI31 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<50> 0 net230
***+  bank16mx1n
***XI27 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<44> 0 net230
***+  bank16mx1n
***XI25 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<63> 0 net230
***+  bank16mx1n
***XI30 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<34> 0 net230
***+  bank16mx1n
***XI19 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<47> 0 net230
***+  bank16mx1n
***XI26 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<61> 0 net230
***+  bank16mx1n
***XI24 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<60> 0 net230
***+  bank16mx1n
***XI34 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<55> 0 net230
***+  bank16mx1n
***XI23 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<48> 0 net230
***+  bank16mx1n
***XI17 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<45> 0 net230
***+  bank16mx1n
***XI3 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<14> 0 net230
***+  bank16mx1n
***XI5 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<13> 0 net230
***+  bank16mx1n
***XI2 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<1> 0 net230
***+  bank16mx1n
***XI1 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<15> 0 net230
***+  bank16mx1n
***XI0 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<0> io_x net230
***+  bank16mx1n
***XI11 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<30> 0 net230
***+  bank16mx1n
***XI10 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<17> 0 net230
***+  bank16mx1n
***XI8 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<16> 0 net230
***+  bank16mx1n
***XI15 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<28> 0 net230
***+  bank16mx1n
***XI9 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<31> 0 net230
***+  bank16mx1n
***XI13 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<29> 0 net230
***+  bank16mx1n
***XI7 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<12> 0 net230
***+  bank16mx1n
***XI6 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<3> 0 net230
***+  bank16mx1n
***XI14 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<19> 0 net230
***+  bank16mx1n
***XI4 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<2> 0 net230
***+  bank16mx1n
***XI12 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<18> 0 net230
***+  bank16mx1n
***XI39 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<56> 0 net230
***+  bank16mx1n
***XI16 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<46> 0 net230
***+  bank16mx1n
***XI37 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<57> 0 net230
***+  bank16mx1n
***XI29 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<51> 0 net230
***+  bank16mx1n
***XI43 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<58> 0 net230
***+  bank16mx1n
***XI45 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<43> 0 net230
***+  bank16mx1n
***XI46 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<37> 0 net230
***+  bank16mx1n
***XI33 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<38> 0 net230
***+  bank16mx1n
***XI44 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<36> 0 net230
***+  bank16mx1n
XI73 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> net230 net474   atd18
XI160 net476 net493   inv Ln=0.35u Wn=20u M=2 Lp=0.35u Wp=40u
XI310 w_ net480   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI309 net480 net230   inv Ln=0.35u Wn=20u M=2 Lp=0.35u Wp=40u
XI83 d net476   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI221 net491 net485   inv Ln=0.35u Wn=7u M=6 Lp=0.35u Wp=14u
XI159 net230 net487   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI222 net485 q   inv Ln=0.35u Wn=7u M=12 Lp=0.35u Wp=14u
XI223 net496 net491   inv Ln=0.35u Wn=7u M=2 Lp=0.35u Wp=14u
XI161 io_x net493 net487 net230   ctg Lp=0.35u Wp=3.5u Ln=0.35u Wn=3.5u
XI74 net500 io_x  net496   dff1
XI72 net501 net500 net503   sen_ena
XI71 net474 net503   xvald
XI68 a<29> a<28> a<27> a<26> a<25> a<24> ena en<63> en<62> en<61> en<60>
+en<59> en<58> en<57> en<56> en<55> en<54> en<53> en<52> en<51> en<50> en<49>
+en<48> en<47> en<46> en<45> en<44> en<43> en<42> en<41> en<40> en<39> en<38>
+en<37> en<36> en<35> en<34> en<33> en<32> en<31> en<30> en<29> en<28> en<27>
+en<26> en<25> en<24> en<23> en<22> en<21> en<20> en<19> en<18> en<17> en<16>
+en<15> en<14> en<13> en<12> en<11> en<10> en<9> en<8> en<7> en<6> en<5> en<4>
+en<3> en<2> en<1> en<0>   decoder6_64
.ENDS
