************************************************************************
* auCdl Netlist:
*
* Library Name: Lassen_DRAMB
* Top Cell Name: dram1gbn
* View Name: schematic
* Netlisted on: Dec 18 16:47:09 2000
************************************************************************


.GLOBAL vddh! gnd! vbb! vdd! vddh2!

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: ctg
* View Name: schematic
************************************************************************

.SUBCKT ctg C1 C2 N P
MM0 C2 N C1 vbb! NMOS W=Wn L=Ln M=1
MM1 C2 P C1 vdd! PMOS W=Wp L=Lp M=1.0
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: inv
* View Name: schematic
************************************************************************

.SUBCKT inv A Y
MM1 Y A vdd! vdd! PMOS W=Wp L=Lp M=M
MM12 Y A gnd! vbb! NMOS W=Wn L=Ln M=M
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: main_sense
* View Name: schematic
************************************************************************

.SUBCKT main_sense ena io io_ o o_ pre
XI165 pre net20   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
MM5 o pre o_ vbb! NMOS W=1.4u L=350.00n M=1
MM2 o_ io net21 vbb! NMOS W=7u L=350.00n M=1
MM3 o io_ net21 vbb! NMOS W=7u L=350.00n M=1
MM4 net21 ena gnd! vbb! NMOS W=7u L=350.00n M=1
MM0 vdd! o_ o vdd! PMOS W=14u L=350.00n M=1
MM1 o_ net20 o vdd! PMOS W=1.4u L=350.00n M=1
MM17 vdd! o o_ vdd! PMOS W=14u L=350.00n M=1
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: precharge
* View Name: schematic
************************************************************************

.SUBCKT precharge bl bl_ pre
MM4 vddh! pre bl vbb! NMOS W=1.4u L=350.00n M=1
MM6 vddh! pre bl_ vbb! NMOS W=1.4u L=350.00n M=1
MM3 bl pre bl_ vbb! NMOS W=1.4u L=350.00n M=1
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: io
* View Name: schematic
************************************************************************

.SUBCKT io a0 i_o io io_ main_ena pre w_
MM0 net52 net107 gnd! vbb! NMOS W=1.4u L=350.00n M=1
MM12 i_o net93 net52 vbb! NMOS W=1.4u L=350.00n M=1
MM1 i_o net101 net63 vdd! PMOS W=3.5u L=350.00n M=1
MM2 net63 net107 vdd! vdd! PMOS W=3.5u L=350.00n M=1
XI210 main_ena io io_ net73 net70 pre   main_sense
XI218 net73 net83 net111 a0   ctg Lp=0.35u Wp=3.5u Ln=0.35u Wn=3.5u
XI196 io_ net95 a0 net119   ctg Lp=0.35u Wp=3.5u Ln=0.35u Wn=3.5u
XI164 io net95 net119 a0   ctg Lp=0.35u Wp=3.5u Ln=0.35u Wn=3.5u
XI161 net95 i_o net101 net93   ctg Lp=0.35u Wp=3.5u Ln=0.35u Wn=3.5u
XI217 net70 net83 a0 net111   ctg Lp=0.35u Wp=3.5u Ln=0.35u Wn=3.5u
XI224 net83 net107   inv Ln=0.35u Wn=1.4u M=1 Lp=0.35u Wp=2.8u
XI306 w_ net101   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI165 a0 net119   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI307 net101 net93   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI219 a0 net111   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI195 io io_ pre   precharge
CC20 io_ gnd! 200f $[CP]
CC22 io gnd! 200f $[CP]
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: nand2
* View Name: schematic
************************************************************************

.SUBCKT nand2 A B Y
MM14 net28 B gnd! vbb! NMOS W=Wn L=Ln M=1
MM13 Y A net28 vbb! NMOS W=Wn L=Ln M=1
MM12 Y A vdd! vdd! PMOS W=Wp L=Lp M=1.0
MM11 Y B vdd! vdd! PMOS W=Wp L=Lp M=1.0
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: nor3
* View Name: schematic
************************************************************************

.SUBCKT nor3 A B C Y
MM16 Y C gnd! vbb! NMOS W=Wn L=Ln M=1
MM17 Y B gnd! vbb! NMOS W=Wn L=Ln M=1
MM18 Y A gnd! vbb! NMOS W=Wn L=Ln M=1
MM9 net29 C vdd! vdd! PMOS W=Wp L=Lp M=1.0
MM10 net25 B net29 vdd! PMOS W=Wp L=Lp M=1.0
MM15 Y A net25 vdd! PMOS W=Wp L=Lp M=1.0
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: nand5
* View Name: schematic
************************************************************************

.SUBCKT nand5 A B C D E Y
MM3 net40 D net12 vbb! NMOS W=Wn L=Ln M=1
MM1 net60 C net40 vbb! NMOS W=Wn L=Ln M=1
MM14 net28 B net60 vbb! NMOS W=Wn L=Ln M=1
MM13 Y A net28 vbb! NMOS W=Wn L=Ln M=1
MM4 net12 E gnd! vbb! NMOS W=Wn L=Ln M=1
MM5 Y E vdd! vdd! PMOS W=Wp L=Lp M=1
MM2 Y D vdd! vdd! PMOS W=Wp L=Lp M=1
MM0 Y C vdd! vdd! PMOS W=Wp L=Lp M=1
MM12 Y A vdd! vdd! PMOS W=Wp L=Lp M=1
MM11 Y B vdd! vdd! PMOS W=Wp L=Lp M=1
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: nor4
* View Name: schematic
************************************************************************

.SUBCKT nor4 A B C D Y
MM19 gnd! A Y vbb! NMOS W=Wn L=Ln M=1
MM18 gnd! B Y vbb! NMOS W=Wn L=Ln M=1
MM17 gnd! C Y vbb! NMOS W=Wn L=Ln M=1
MM16 gnd! D Y vbb! NMOS W=Wn L=Ln M=1
MM8 vdd! D net35 vdd! PMOS W=Wp L=Lp M=1.0
MM9 net35 C net31 vdd! PMOS W=Wp L=Lp M=1.0
MM15 net27 A Y vdd! PMOS W=Wp L=Lp M=1.0
MM10 net31 B net27 vdd! PMOS W=Wp L=Lp M=1.0
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: delay10
* View Name: schematic
************************************************************************

.SUBCKT delay10 A Y
XI47 net011 net39   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI57 net017 Y   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI45 net39 net40   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI44 net40 net023   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI48 net023 net04   inv Ln=2.5u Wn=1u M=1 Lp=2.5u Wp=1u
XI51 net04 net12   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI52 net9 net029   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI53 net029 net017   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI46 A net011   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI50 net12 net9   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: atd1
* View Name: schematic
************************************************************************

.SUBCKT atd1 A Y
XI58 net32 net22   delay10
XI59 net38 net24   delay10
MM1 net38 net22 net39 vbb! NMOS W=1.4u L=350.00n M=1
MM0 net39 net24 net32 vbb! NMOS W=1.4u L=350.00n M=1
XI68 A net32   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI62 net20 Y   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI69 net39 net20   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI46 net32 net38   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
.ENDS

************************************************************************
* Library Name: Lassen_DRAMB
* Cell Name: atd18m
* View Name: schematic
************************************************************************

.SUBCKT atd18m a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7>
+a<6> a<5> a<4> a<3> a<2> a<1> a<0> ena w_ y
XI75 net137 ena net159   nand2 Lp=0.35u Wp=16u Ln=0.35u Wn=8u
XI103 net99 net97 net189 net163   nor3 Lp=0.35u Wp=7u Ln=0.35u Wn=3.5u
XI74 net157 net152 net147 net142 net163 net137   nand5 Lp=0.35u Wp=4u Ln=0.35u
+Wn=7u
XI96 net169 net165 net171 net167 net142   nor4 Lp=0.35u Wp=7u Ln=0.35u Wn=3.5u
XI93 net181 net183 net187 net185 net152   nor4 Lp=0.35u Wp=7u Ln=0.35u Wn=3.5u
XI92 net193 net195 net197 net191 net157   nor4 Lp=0.35u Wp=7u Ln=0.35u Wn=3.5u
XI94 net175 net179 net173 net177 net147   nor4 Lp=0.35u Wp=7u Ln=0.35u Wn=3.5u
XI81 net159 y   inv Ln=0.35u Wn=8u M=9 Lp=0.35u Wp=16u
XI101 a<16> net99   atd1
XI102 a<17> net97   atd1
XI97 a<14> net171   atd1
XI98 a<12> net169   atd1
XI71 a<3> net191   atd1
XI99 a<15> net167   atd1
XI79 w_ net189   atd1
XI91 a<10> net173   atd1
XI68 a<0> net193   atd1
XI83 a<4> net181   atd1
XI84 a<5> net183   atd1
XI82 a<7> net185   atd1
XI88 a<8> net175   atd1
XI85 a<6> net187   atd1
XI100 a<13> net165   atd1
XI69 a<1> net195   atd1
XI70 a<2> net197   atd1
XI90 a<11> net177   atd1
XI89 a<9> net179   atd1
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: col_sel1m
* View Name: schematic
************************************************************************

.SUBCKT col_sel1m a0 a1 a2 ena pre wl xvld
c1 pre 0 1pf
XI32 a0 a1 a2 xvld ena net119  nand5 Lp=0.35u Wp=4u Ln=0.35u Wn=10u
MM17 wl net119 gnd! vbb! NMOS W=14u L=350.00n M=1
MM8  wl net119 vddh2! vddh2! PMOS W=28u L=350.00n M=1.0
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: col_sel3_8m
* View Name: schematic
************************************************************************

.SUBCKT col_sel3_8m a<2> a<1> a<0> cs<7> cs<6> cs<5> cs<4> cs<3> cs<2> cs<1>
+cs<0> ena pre xvld
XI51 net33 net31 net25 ena pre cs<7> xvld   col_sel1m
XI41 net35 net29 net27 ena pre cs<0> xvld   col_sel1m
XI49 net35 net31 net27 ena pre cs<2> xvld   col_sel1m
XI50 net35 net31 net25 ena pre cs<6> xvld   col_sel1m
XI47 net33 net29 net27 ena pre cs<1> xvld   col_sel1m
XI52 net33 net29 net25 ena pre cs<5> xvld   col_sel1m
XI48 net33 net31 net27 ena pre cs<3> xvld   col_sel1m
XI53 net35 net29 net25 ena pre cs<4> xvld   col_sel1m
XI88 net35 net33   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI56 a<2> net27   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI90 a<0> net35   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI57 net27 net25   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI54 net29 net31   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI55 a<1> net29   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: decoder4_16
* View Name: schematic
************************************************************************

.SUBCKT decoder4_16 A<3> A<2> A<1> A<0> ENA X<15> X<14> X<13> X<12> X<11>
+X<10> X<9> X<8> X<7> X<6> X<5> X<4> X<3> X<2> X<1> X<0>
XI27 net146 net142 net138 net132 net128 net126   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI17 net146 net117 net138 net134 net128 net131   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI32 net146 net142 net136 net132 net130 net286   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI31 net146 net142 net136 net132 net128 net285   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI30 net146 net142 net136 net134 net130 net150   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI29 net146 net142 net136 net134 net128 net156   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI23 net146 net117 net136 net132 net128 net162   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI19 net146 net117 net138 net132 net128 net168   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI24 net146 net117 net136 net132 net130 net174   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI20 net146 net117 net138 net132 net130 net180   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI21 net146 net117 net136 net134 net128 net186   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI22 net146 net117 net136 net134 net130 net192   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI18 net146 net117 net138 net134 net130 net198   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI26 net146 net142 net138 net134 net130 net204   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI28 net146 net142 net138 net132 net130 net210   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI25 net146 net142 net138 net134 net128 net216   nand5 Lp=0.35u Wp=2.1u
+Ln=0.35u Wn=2.1u
XI93 ENA net144   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=4.2u
XI45 net198 X<14>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI46 net168 X<13>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI47 net180 X<12>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI44 net131 X<15>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI48 net186 X<11>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI49 net192 X<10>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI50 net162 X<9>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI51 net174 X<8>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI52 net216 X<7>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI53 net204 X<6>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI54 net126 X<5>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI55 net210 X<4>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI56 net156 X<3>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI57 net150 X<2>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI58 net285 X<1>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI59 net286 X<0>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI42 net144 net146   inv Ln=0.35u Wn=2.1u M=3 Lp=0.35u Wp=4.2u
XI41 A<1> net132   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=3.2u
XI40 net132 net134   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=3.2u
XI39 net130 net128   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=3.2u
XI38 A<0> net130   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=3.2u
XI37 A<2> net136   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=3.2u
XI33 A<3> net142   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=3.2u
XI36 net136 net138   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=3.2u
XI35 net142 net117   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=3.2u
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: col_sel7_128
* View Name: schematic
************************************************************************

.SUBCKT col_sel7_128 a<6> a<5> a<4> a<3> a<2> a<1> a<0> cs<127> cs<126>
+cs<125> cs<124> cs<123> cs<122> cs<121> cs<120> cs<119> cs<118> cs<117>
+cs<116> cs<115> cs<114> cs<113> cs<112> cs<111> cs<110> cs<109> cs<108>
+cs<107> cs<106> cs<105> cs<104> cs<103> cs<102> cs<101> cs<100> cs<99> cs<98>
+cs<97> cs<96> cs<95> cs<94> cs<93> cs<92> cs<91> cs<90> cs<89> cs<88> cs<87>
+cs<86> cs<85> cs<84> cs<83> cs<82> cs<81> cs<80> cs<79> cs<78> cs<77> cs<76>
+cs<75> cs<74> cs<73> cs<72> cs<71> cs<70> cs<69> cs<68> cs<67> cs<66> cs<65>
+cs<64> cs<63> cs<62> cs<61> cs<60> cs<59> cs<58> cs<57> cs<56> cs<55> cs<54>
+cs<53> cs<52> cs<51> cs<50> cs<49> cs<48> cs<47> cs<46> cs<45> cs<44> cs<43>
+cs<42> cs<41> cs<40> cs<39> cs<38> cs<37> cs<36> cs<35> cs<34> cs<33> cs<32>
+cs<31> cs<30> cs<29> cs<28> cs<27> cs<26> cs<25> cs<24> cs<23> cs<22> cs<21>
+cs<20> cs<19> cs<18> cs<17> cs<16> cs<15> cs<14> cs<13> cs<12> cs<11> cs<10>
+cs<9> cs<8> cs<7> cs<6> cs<5> cs<4> cs<3> cs<2> cs<1> cs<0> ena pre xvld
XI72 a<2> a<1> a<0> cs<127> cs<126> cs<125> cs<124> cs<123> cs<122> cs<121>
+cs<120> net<15> net201 net213   col_sel3_8m
XI73 a<2> a<1> a<0> cs<95> cs<94> cs<93> cs<92> cs<91> cs<90> cs<89> cs<88>
+net<11> net201 net213   col_sel3_8m
XI74 a<2> a<1> a<0> cs<87> cs<86> cs<85> cs<84> cs<83> cs<82> cs<81> cs<80>
+net<10> net201 net213   col_sel3_8m
XI75 a<2> a<1> a<0> cs<79> cs<78> cs<77> cs<76> cs<75> cs<74> cs<73> cs<72>
+net<9> net201 net213   col_sel3_8m
XI76 a<2> a<1> a<0> cs<103> cs<102> cs<101> cs<100> cs<99> cs<98> cs<97>
+cs<96> net<12> net201 net213   col_sel3_8m
XI77 a<2> a<1> a<0> cs<119> cs<118> cs<117> cs<116> cs<115> cs<114> cs<113>
+cs<112> net<14> net201 net213   col_sel3_8m
XI78 a<2> a<1> a<0> cs<111> cs<110> cs<109> cs<108> cs<107> cs<106> cs<105>
+cs<104> net<13> net201 net213   col_sel3_8m
XI71 a<2> a<1> a<0> cs<71> cs<70> cs<69> cs<68> cs<67> cs<66> cs<65> cs<64>
+net<8> net201 net213   col_sel3_8m
XI63 a<2> a<1> a<0> cs<7> cs<6> cs<5> cs<4> cs<3> cs<2> cs<1> cs<0> net<0>
+net110 net108   col_sel3_8m
XI70 a<2> a<1> a<0> cs<63> cs<62> cs<61> cs<60> cs<59> cs<58> cs<57> cs<56>
+net<7> net110 net108   col_sel3_8m
XI66 a<2> a<1> a<0> cs<31> cs<30> cs<29> cs<28> cs<27> cs<26> cs<25> cs<24>
+net<3> net110 net108   col_sel3_8m
XI65 a<2> a<1> a<0> cs<23> cs<22> cs<21> cs<20> cs<19> cs<18> cs<17> cs<16>
+net<2> net110 net108   col_sel3_8m
XI64 a<2> a<1> a<0> cs<15> cs<14> cs<13> cs<12> cs<11> cs<10> cs<9> cs<8>
+net<1> net110 net108   col_sel3_8m
XI67 a<2> a<1> a<0> cs<39> cs<38> cs<37> cs<36> cs<35> cs<34> cs<33> cs<32>
+net<4> net110 net108   col_sel3_8m
XI69 a<2> a<1> a<0> cs<55> cs<54> cs<53> cs<52> cs<51> cs<50> cs<49> cs<48>
+net<6> net110 net108   col_sel3_8m
XI68 a<2> a<1> a<0> cs<47> cs<46> cs<45> cs<44> cs<43> cs<42> cs<41> cs<40>
+net<5> net110 net108   col_sel3_8m
XI61 a<6> a<5> a<4> a<3> ena net<15> net<14> net<13> net<12> net<11> net<10>
+net<9> net<8> net<7> net<6> net<5> net<4> net<3> net<2> net<1> net<0>  
+decoder4_16
XI81 pre net199   inv Ln=0.35u Wn=8u M=27 Lp=0.35u Wp=16u
XI84 xvld net211   inv Ln=0.35u Wn=10u M=6 Lp=0.35u Wp=20u
XI55 pre net112   inv Ln=0.35u Wn=8u M=27 Lp=0.35u Wp=16u
XI54 net112 net110   inv Ln=0.35u Wn=8u M=81 Lp=0.35u Wp=16u
XI82 net199 net201   inv Ln=0.35u Wn=8u M=81 Lp=0.35u Wp=16u
XI79 net106 net108   inv Ln=0.35u Wn=10u M=18 Lp=0.35u Wp=20u
XI80 xvld net106   inv Ln=0.35u Wn=10u M=6 Lp=0.35u Wp=20u
XI83 net211 net213   inv Ln=0.35u Wn=10u M=18 Lp=0.35u Wp=20u
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: nand3
* View Name: schematic
************************************************************************

.SUBCKT nand3 A B C Y
MM1 net60 C gnd! vbb! NMOS W=Wn L=Ln M=1
MM14 net28 B net60 vbb! NMOS W=Wn L=Ln M=1
MM13 Y A net28 vbb! NMOS W=Wn L=Ln M=1
MM0 Y C vdd! vdd! PMOS W=Wp L=Lp M=1.0
MM12 Y A vdd! vdd! PMOS W=Wp L=Lp M=1.0
MM11 Y B vdd! vdd! PMOS W=Wp L=Lp M=1.0
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: decoder2_4
* View Name: schematic
************************************************************************

.SUBCKT decoder2_4 A<1> A<0> ENA X<3> X<2> X<1> X<0>
XI32 net132 net142 net136 net286   nand3 Lp=0.35u Wp=2.1u Ln=0.35u Wn=2.1u
XI31 net132 net128 net136 net285   nand3 Lp=0.35u Wp=2.1u Ln=0.35u Wn=2.1u
XI30 net134 net142 net136 net150   nand3 Lp=0.35u Wp=2.1u Ln=0.35u Wn=2.1u
XI29 net134 net128 net136 net156   nand3 Lp=0.35u Wp=2.1u Ln=0.35u Wn=2.1u
XI93 ENA net144   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=4.2u
XI56 net156 X<3>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI57 net150 X<2>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI58 net285 X<1>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI59 net286 X<0>   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI42 net144 net136   inv Ln=0.35u Wn=2.1u M=3 Lp=0.35u Wp=4.2u
XI41 A<1> net132   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=3.2u
XI40 net132 net134   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=3.2u
XI39 net142 net128   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=3.2u
XI38 A<0> net142   inv Ln=0.35u Wn=2.1u M=1 Lp=0.35u Wp=3.2u
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: col_sel9_512
* View Name: schematic
************************************************************************

.SUBCKT col_sel9_512 a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> cs<511>
+cs<510> cs<509> cs<508> cs<507> cs<506> cs<505> cs<504> cs<503> cs<502>
+cs<501> cs<500> cs<499> cs<498> cs<497> cs<496> cs<495> cs<494> cs<493>
+cs<492> cs<491> cs<490> cs<489> cs<488> cs<487> cs<486> cs<485> cs<484>
+cs<483> cs<482> cs<481> cs<480> cs<479> cs<478> cs<477> cs<476> cs<475>
+cs<474> cs<473> cs<472> cs<471> cs<470> cs<469> cs<468> cs<467> cs<466>
+cs<465> cs<464> cs<463> cs<462> cs<461> cs<460> cs<459> cs<458> cs<457>
+cs<456> cs<455> cs<454> cs<453> cs<452> cs<451> cs<450> cs<449> cs<448>
+cs<447> cs<446> cs<445> cs<444> cs<443> cs<442> cs<441> cs<440> cs<439>
+cs<438> cs<437> cs<436> cs<435> cs<434> cs<433> cs<432> cs<431> cs<430>
+cs<429> cs<428> cs<427> cs<426> cs<425> cs<424> cs<423> cs<422> cs<421>
+cs<420> cs<419> cs<418> cs<417> cs<416> cs<415> cs<414> cs<413> cs<412>
+cs<411> cs<410> cs<409> cs<408> cs<407> cs<406> cs<405> cs<404> cs<403>
+cs<402> cs<401> cs<400> cs<399> cs<398> cs<397> cs<396> cs<395> cs<394>
+cs<393> cs<392> cs<391> cs<390> cs<389> cs<388> cs<387> cs<386> cs<385>
+cs<384> cs<383> cs<382> cs<381> cs<380> cs<379> cs<378> cs<377> cs<376>
+cs<375> cs<374> cs<373> cs<372> cs<371> cs<370> cs<369> cs<368> cs<367>
+cs<366> cs<365> cs<364> cs<363> cs<362> cs<361> cs<360> cs<359> cs<358>
+cs<357> cs<356> cs<355> cs<354> cs<353> cs<352> cs<351> cs<350> cs<349>
+cs<348> cs<347> cs<346> cs<345> cs<344> cs<343> cs<342> cs<341> cs<340>
+cs<339> cs<338> cs<337> cs<336> cs<335> cs<334> cs<333> cs<332> cs<331>
+cs<330> cs<329> cs<328> cs<327> cs<326> cs<325> cs<324> cs<323> cs<322>
+cs<321> cs<320> cs<319> cs<318> cs<317> cs<316> cs<315> cs<314> cs<313>
+cs<312> cs<311> cs<310> cs<309> cs<308> cs<307> cs<306> cs<305> cs<304>
+cs<303> cs<302> cs<301> cs<300> cs<299> cs<298> cs<297> cs<296> cs<295>
+cs<294> cs<293> cs<292> cs<291> cs<290> cs<289> cs<288> cs<287> cs<286>
+cs<285> cs<284> cs<283> cs<282> cs<281> cs<280> cs<279> cs<278> cs<277>
+cs<276> cs<275> cs<274> cs<273> cs<272> cs<271> cs<270> cs<269> cs<268>
+cs<267> cs<266> cs<265> cs<264> cs<263> cs<262> cs<261> cs<260> cs<259>
+cs<258> cs<257> cs<256> cs<255> cs<254> cs<253> cs<252> cs<251> cs<250>
+cs<249> cs<248> cs<247> cs<246> cs<245> cs<244> cs<243> cs<242> cs<241>
+cs<240> cs<239> cs<238> cs<237> cs<236> cs<235> cs<234> cs<233> cs<232>
+cs<231> cs<230> cs<229> cs<228> cs<227> cs<226> cs<225> cs<224> cs<223>
+cs<222> cs<221> cs<220> cs<219> cs<218> cs<217> cs<216> cs<215> cs<214>
+cs<213> cs<212> cs<211> cs<210> cs<209> cs<208> cs<207> cs<206> cs<205>
+cs<204> cs<203> cs<202> cs<201> cs<200> cs<199> cs<198> cs<197> cs<196>
+cs<195> cs<194> cs<193> cs<192> cs<191> cs<190> cs<189> cs<188> cs<187>
+cs<186> cs<185> cs<184> cs<183> cs<182> cs<181> cs<180> cs<179> cs<178>
+cs<177> cs<176> cs<175> cs<174> cs<173> cs<172> cs<171> cs<170> cs<169>
+cs<168> cs<167> cs<166> cs<165> cs<164> cs<163> cs<162> cs<161> cs<160>
+cs<159> cs<158> cs<157> cs<156> cs<155> cs<154> cs<153> cs<152> cs<151>
+cs<150> cs<149> cs<148> cs<147> cs<146> cs<145> cs<144> cs<143> cs<142>
+cs<141> cs<140> cs<139> cs<138> cs<137> cs<136> cs<135> cs<134> cs<133>
+cs<132> cs<131> cs<130> cs<129> cs<128> cs<127> cs<126> cs<125> cs<124>
+cs<123> cs<122> cs<121> cs<120> cs<119> cs<118> cs<117> cs<116> cs<115>
+cs<114> cs<113> cs<112> cs<111> cs<110> cs<109> cs<108> cs<107> cs<106>
+cs<105> cs<104> cs<103> cs<102> cs<101> cs<100> cs<99> cs<98> cs<97> cs<96>
+cs<95> cs<94> cs<93> cs<92> cs<91> cs<90> cs<89> cs<88> cs<87> cs<86> cs<85>
+cs<84> cs<83> cs<82> cs<81> cs<80> cs<79> cs<78> cs<77> cs<76> cs<75> cs<74>
+cs<73> cs<72> cs<71> cs<70> cs<69> cs<68> cs<67> cs<66> cs<65> cs<64> cs<63>
+cs<62> cs<61> cs<60> cs<59> cs<58> cs<57> cs<56> cs<55> cs<54> cs<53> cs<52>
+cs<51> cs<50> cs<49> cs<48> cs<47> cs<46> cs<45> cs<44> cs<43> cs<42> cs<41>
+cs<40> cs<39> cs<38> cs<37> cs<36> cs<35> cs<34> cs<33> cs<32> cs<31> cs<30>
+cs<29> cs<28> cs<27> cs<26> cs<25> cs<24> cs<23> cs<22> cs<21> cs<20> cs<19>
+cs<18> cs<17> cs<16> cs<15> cs<14> cs<13> cs<12> cs<11> cs<10> cs<9> cs<8>
+cs<7> cs<6> cs<5> cs<4> cs<3> cs<2> cs<1> cs<0> ena pre xvld
XI63 a<6> a<5> a<4> a<3> a<2> a<1> a<0> cs<127> cs<126> cs<125> cs<124>
+cs<123> cs<122> cs<121> cs<120> cs<119> cs<118> cs<117> cs<116> cs<115>
+cs<114> cs<113> cs<112> cs<111> cs<110> cs<109> cs<108> cs<107> cs<106>
+cs<105> cs<104> cs<103> cs<102> cs<101> cs<100> cs<99> cs<98> cs<97> cs<96>
+cs<95> cs<94> cs<93> cs<92> cs<91> cs<90> cs<89> cs<88> cs<87> cs<86> cs<85>
+cs<84> cs<83> cs<82> cs<81> cs<80> cs<79> cs<78> cs<77> cs<76> cs<75> cs<74>
+cs<73> cs<72> cs<71> cs<70> cs<69> cs<68> cs<67> cs<66> cs<65> cs<64> cs<63>
+cs<62> cs<61> cs<60> cs<59> cs<58> cs<57> cs<56> cs<55> cs<54> cs<53> cs<52>
+cs<51> cs<50> cs<49> cs<48> cs<47> cs<46> cs<45> cs<44> cs<43> cs<42> cs<41>
+cs<40> cs<39> cs<38> cs<37> cs<36> cs<35> cs<34> cs<33> cs<32> cs<31> cs<30>
+cs<29> cs<28> cs<27> cs<26> cs<25> cs<24> cs<23> cs<22> cs<21> cs<20> cs<19>
+cs<18> cs<17> cs<16> cs<15> cs<14> cs<13> cs<12> cs<11> cs<10> cs<9> cs<8>
+cs<7> cs<6> cs<5> cs<4> cs<3> cs<2> cs<1> cs<0> net<0> net110 net108  
+col_sel7_128
XI66 a<6> a<5> a<4> a<3> a<2> a<1> a<0> cs<511> cs<510> cs<509> cs<508>
+cs<507> cs<506> cs<505> cs<504> cs<503> cs<502> cs<501> cs<500> cs<499>
+cs<498> cs<497> cs<496> cs<495> cs<494> cs<493> cs<492> cs<491> cs<490>
+cs<489> cs<488> cs<487> cs<486> cs<485> cs<484> cs<483> cs<482> cs<481>
+cs<480> cs<479> cs<478> cs<477> cs<476> cs<475> cs<474> cs<473> cs<472>
+cs<471> cs<470> cs<469> cs<468> cs<467> cs<466> cs<465> cs<464> cs<463>
+cs<462> cs<461> cs<460> cs<459> cs<458> cs<457> cs<456> cs<455> cs<454>
+cs<453> cs<452> cs<451> cs<450> cs<449> cs<448> cs<447> cs<446> cs<445>
+cs<444> cs<443> cs<442> cs<441> cs<440> cs<439> cs<438> cs<437> cs<436>
+cs<435> cs<434> cs<433> cs<432> cs<431> cs<430> cs<429> cs<428> cs<427>
+cs<426> cs<425> cs<424> cs<423> cs<422> cs<421> cs<420> cs<419> cs<418>
+cs<417> cs<416> cs<415> cs<414> cs<413> cs<412> cs<411> cs<410> cs<409>
+cs<408> cs<407> cs<406> cs<405> cs<404> cs<403> cs<402> cs<401> cs<400>
+cs<399> cs<398> cs<397> cs<396> cs<395> cs<394> cs<393> cs<392> cs<391>
+cs<390> cs<389> cs<388> cs<387> cs<386> cs<385> cs<384> net<3> net110 net108
+  col_sel7_128
XI65 a<6> a<5> a<4> a<3> a<2> a<1> a<0> cs<383> cs<382> cs<381> cs<380>
+cs<379> cs<378> cs<377> cs<376> cs<375> cs<374> cs<373> cs<372> cs<371>
+cs<370> cs<369> cs<368> cs<367> cs<366> cs<365> cs<364> cs<363> cs<362>
+cs<361> cs<360> cs<359> cs<358> cs<357> cs<356> cs<355> cs<354> cs<353>
+cs<352> cs<351> cs<350> cs<349> cs<348> cs<347> cs<346> cs<345> cs<344>
+cs<343> cs<342> cs<341> cs<340> cs<339> cs<338> cs<337> cs<336> cs<335>
+cs<334> cs<333> cs<332> cs<331> cs<330> cs<329> cs<328> cs<327> cs<326>
+cs<325> cs<324> cs<323> cs<322> cs<321> cs<320> cs<319> cs<318> cs<317>
+cs<316> cs<315> cs<314> cs<313> cs<312> cs<311> cs<310> cs<309> cs<308>
+cs<307> cs<306> cs<305> cs<304> cs<303> cs<302> cs<301> cs<300> cs<299>
+cs<298> cs<297> cs<296> cs<295> cs<294> cs<293> cs<292> cs<291> cs<290>
+cs<289> cs<288> cs<287> cs<286> cs<285> cs<284> cs<283> cs<282> cs<281>
+cs<280> cs<279> cs<278> cs<277> cs<276> cs<275> cs<274> cs<273> cs<272>
+cs<271> cs<270> cs<269> cs<268> cs<267> cs<266> cs<265> cs<264> cs<263>
+cs<262> cs<261> cs<260> cs<259> cs<258> cs<257> cs<256> net<2> net110 net108
+  col_sel7_128
XI64 a<6> a<5> a<4> a<3> a<2> a<1> a<0> cs<255> cs<254> cs<253> cs<252>
+cs<251> cs<250> cs<249> cs<248> cs<247> cs<246> cs<245> cs<244> cs<243>
+cs<242> cs<241> cs<240> cs<239> cs<238> cs<237> cs<236> cs<235> cs<234>
+cs<233> cs<232> cs<231> cs<230> cs<229> cs<228> cs<227> cs<226> cs<225>
+cs<224> cs<223> cs<222> cs<221> cs<220> cs<219> cs<218> cs<217> cs<216>
+cs<215> cs<214> cs<213> cs<212> cs<211> cs<210> cs<209> cs<208> cs<207>
+cs<206> cs<205> cs<204> cs<203> cs<202> cs<201> cs<200> cs<199> cs<198>
+cs<197> cs<196> cs<195> cs<194> cs<193> cs<192> cs<191> cs<190> cs<189>
+cs<188> cs<187> cs<186> cs<185> cs<184> cs<183> cs<182> cs<181> cs<180>
+cs<179> cs<178> cs<177> cs<176> cs<175> cs<174> cs<173> cs<172> cs<171>
+cs<170> cs<169> cs<168> cs<167> cs<166> cs<165> cs<164> cs<163> cs<162>
+cs<161> cs<160> cs<159> cs<158> cs<157> cs<156> cs<155> cs<154> cs<153>
+cs<152> cs<151> cs<150> cs<149> cs<148> cs<147> cs<146> cs<145> cs<144>
+cs<143> cs<142> cs<141> cs<140> cs<139> cs<138> cs<137> cs<136> cs<135>
+cs<134> cs<133> cs<132> cs<131> cs<130> cs<129> cs<128> net<1> net110 net108
+  col_sel7_128
XI61 a<8> a<7> ena net<3> net<2> net<1> net<0>   decoder2_4
XI55 pre net112   inv Ln=0.35u Wn=8u M=9 Lp=0.35u Wp=16u
XI54 net112 net110   inv Ln=0.35u Wn=8u M=27 Lp=0.35u Wp=16u
XI79 net106 net108   inv Ln=0.35u Wn=8u M=6 Lp=0.35u Wp=16u
XI80 xvld net106   inv Ln=0.35u Wn=10u M=2 Lp=0.35u Wp=20u
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: deco1m
* View Name: schematic
************************************************************************

.SUBCKT deco1m a0 a1 a2 ena pre wl xvld
c1 pre 0 1pf
XI32 a0 a1 a2 xvld ena net119  nand5 Lp=0.35u Wp=4u Ln=0.35u Wn=10u
MM17 wl net119 gnd! vbb! NMOS W=14u L=350.00n M=1
MM8  wl net119 vddh2! vddh2! PMOS W=28u L=350.00n M=1.0
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: deco3_8m
* View Name: schematic
************************************************************************

.SUBCKT deco3_8m a<2> a<1> a<0> ena pre wl<7> wl<6> wl<5> wl<4> wl<3> wl<2>
+wl<1> wl<0> xvld
XI51 net33 net31 net25 ena pre wl<7> xvld   deco1m
XI41 net35 net29 net27 ena pre wl<0> xvld   deco1m
XI49 net35 net31 net27 ena pre wl<2> xvld   deco1m
XI50 net35 net31 net25 ena pre wl<6> xvld   deco1m
XI47 net33 net29 net27 ena pre wl<1> xvld   deco1m
XI52 net33 net29 net25 ena pre wl<5> xvld   deco1m
XI48 net33 net31 net27 ena pre wl<3> xvld   deco1m
XI53 net35 net29 net25 ena pre wl<4> xvld   deco1m
XI88 net35 net33   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI56 a<2> net27   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI90 a<0> net35   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI57 net27 net25   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI54 net29 net31   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI55 a<1> net29   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: deco7_128
* View Name: schematic
************************************************************************

.SUBCKT deco7_128 a<6> a<5> a<4> a<3> a<2> a<1> a<0> ena pre wl<127> wl<126>
+wl<125> wl<124> wl<123> wl<122> wl<121> wl<120> wl<119> wl<118> wl<117>
+wl<116> wl<115> wl<114> wl<113> wl<112> wl<111> wl<110> wl<109> wl<108>
+wl<107> wl<106> wl<105> wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98>
+wl<97> wl<96> wl<95> wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87>
+wl<86> wl<85> wl<84> wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76>
+wl<75> wl<74> wl<73> wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65>
+wl<64> wl<63> wl<62> wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54>
+wl<53> wl<52> wl<51> wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43>
+wl<42> wl<41> wl<40> wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32>
+wl<31> wl<30> wl<29> wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21>
+wl<20> wl<19> wl<18> wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10>
+wl<9> wl<8> wl<7> wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0> xvld
XI61 a<6> a<5> a<4> a<3> ena net<15> net<14> net<13> net<12> net<11> net<10>
+net<9> net<8> net<7> net<6> net<5> net<4> net<3> net<2> net<1> net<0>  
+decoder4_16
XI81 pre net199   inv Ln=0.35u Wn=8u M=27 Lp=0.35u Wp=16u
XI84 xvld net211   inv Ln=0.35u Wn=10u M=6 Lp=0.35u Wp=20u
XI55 pre net112   inv Ln=0.35u Wn=8u M=27 Lp=0.35u Wp=16u
XI54 net112 net110   inv Ln=0.35u Wn=8u M=81 Lp=0.35u Wp=16u
XI82 net199 net201   inv Ln=0.35u Wn=8u M=81 Lp=0.35u Wp=16u
XI79 net106 net108   inv Ln=0.35u Wn=10u M=18 Lp=0.35u Wp=20u
XI80 xvld net106   inv Ln=0.35u Wn=10u M=6 Lp=0.35u Wp=20u
XI83 net211 net213   inv Ln=0.35u Wn=10u M=18 Lp=0.35u Wp=20u
XI72 a<2> a<1> a<0> net<15> net201 wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> net213   deco3_8m
XI73 a<2> a<1> a<0> net<11> net201 wl<95> wl<94> wl<93> wl<92> wl<91> wl<90>
+wl<89> wl<88> net213   deco3_8m
XI74 a<2> a<1> a<0> net<10> net201 wl<87> wl<86> wl<85> wl<84> wl<83> wl<82>
+wl<81> wl<80> net213   deco3_8m
XI75 a<2> a<1> a<0> net<9> net201 wl<79> wl<78> wl<77> wl<76> wl<75> wl<74>
+wl<73> wl<72> net213   deco3_8m
XI76 a<2> a<1> a<0> net<12> net201 wl<103> wl<102> wl<101> wl<100> wl<99>
+wl<98> wl<97> wl<96> net213   deco3_8m
XI77 a<2> a<1> a<0> net<14> net201 wl<119> wl<118> wl<117> wl<116> wl<115>
+wl<114> wl<113> wl<112> net213   deco3_8m
XI78 a<2> a<1> a<0> net<13> net201 wl<111> wl<110> wl<109> wl<108> wl<107>
+wl<106> wl<105> wl<104> net213   deco3_8m
XI71 a<2> a<1> a<0> net<8> net201 wl<71> wl<70> wl<69> wl<68> wl<67> wl<66>
+wl<65> wl<64> net213   deco3_8m
XI63 a<2> a<1> a<0> net<0> net110 wl<7> wl<6> wl<5> wl<4> wl<3> wl<2> wl<1>
+wl<0> net108   deco3_8m
XI70 a<2> a<1> a<0> net<7> net110 wl<63> wl<62> wl<61> wl<60> wl<59> wl<58>
+wl<57> wl<56> net108   deco3_8m
XI66 a<2> a<1> a<0> net<3> net110 wl<31> wl<30> wl<29> wl<28> wl<27> wl<26>
+wl<25> wl<24> net108   deco3_8m
XI65 a<2> a<1> a<0> net<2> net110 wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> net108   deco3_8m
XI64 a<2> a<1> a<0> net<1> net110 wl<15> wl<14> wl<13> wl<12> wl<11> wl<10>
+wl<9> wl<8> net108   deco3_8m
XI67 a<2> a<1> a<0> net<4> net110 wl<39> wl<38> wl<37> wl<36> wl<35> wl<34>
+wl<33> wl<32> net108   deco3_8m
XI69 a<2> a<1> a<0> net<6> net110 wl<55> wl<54> wl<53> wl<52> wl<51> wl<50>
+wl<49> wl<48> net108   deco3_8m
XI68 a<2> a<1> a<0> net<5> net110 wl<47> wl<46> wl<45> wl<44> wl<43> wl<42>
+wl<41> wl<40> net108   deco3_8m
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: deco9_512
* View Name: schematic
************************************************************************

.SUBCKT deco9_512 a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> ena pre wl<511>
+wl<510> wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502>
+wl<501> wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493>
+wl<492> wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484>
+wl<483> wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475>
+wl<474> wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466>
+wl<465> wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457>
+wl<456> wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448>
+wl<447> wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439>
+wl<438> wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430>
+wl<429> wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421>
+wl<420> wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412>
+wl<411> wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403>
+wl<402> wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394>
+wl<393> wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385>
+wl<384> wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376>
+wl<375> wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367>
+wl<366> wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358>
+wl<357> wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349>
+wl<348> wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340>
+wl<339> wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331>
+wl<330> wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322>
+wl<321> wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313>
+wl<312> wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304>
+wl<303> wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295>
+wl<294> wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286>
+wl<285> wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277>
+wl<276> wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268>
+wl<267> wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259>
+wl<258> wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250>
+wl<249> wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241>
+wl<240> wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232>
+wl<231> wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223>
+wl<222> wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214>
+wl<213> wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205>
+wl<204> wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196>
+wl<195> wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187>
+wl<186> wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178>
+wl<177> wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169>
+wl<168> wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160>
+wl<159> wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151>
+wl<150> wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142>
+wl<141> wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133>
+wl<132> wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124>
+wl<123> wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115>
+wl<114> wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106>
+wl<105> wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96>
+wl<95> wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85>
+wl<84> wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74>
+wl<73> wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63>
+wl<62> wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52>
+wl<51> wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41>
+wl<40> wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30>
+wl<29> wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19>
+wl<18> wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8>
+wl<7> wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0> xvld
XI61 a<8> a<7> ena net<3> net<2> net<1> net<0>   decoder2_4
XI63 a<6> a<5> a<4> a<3> a<2> a<1> a<0> net<0> net110 wl<127> wl<126> wl<125>
+wl<124> wl<123> wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116>
+wl<115> wl<114> wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107>
+wl<106> wl<105> wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97>
+wl<96> wl<95> wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86>
+wl<85> wl<84> wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75>
+wl<74> wl<73> wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64>
+wl<63> wl<62> wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53>
+wl<52> wl<51> wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42>
+wl<41> wl<40> wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31>
+wl<30> wl<29> wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20>
+wl<19> wl<18> wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9>
+wl<8> wl<7> wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0> net108   deco7_128
XI66 a<6> a<5> a<4> a<3> a<2> a<1> a<0> net<3> net110 wl<511> wl<510> wl<509>
+wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501> wl<500>
+wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492> wl<491>
+wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483> wl<482>
+wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474> wl<473>
+wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465> wl<464>
+wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456> wl<455>
+wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447> wl<446>
+wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438> wl<437>
+wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429> wl<428>
+wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420> wl<419>
+wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411> wl<410>
+wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402> wl<401>
+wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393> wl<392>
+wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384> net108  
+deco7_128
XI65 a<6> a<5> a<4> a<3> a<2> a<1> a<0> net<2> net110 wl<383> wl<382> wl<381>
+wl<380> wl<379> wl<378> wl<377> wl<376> wl<375> wl<374> wl<373> wl<372>
+wl<371> wl<370> wl<369> wl<368> wl<367> wl<366> wl<365> wl<364> wl<363>
+wl<362> wl<361> wl<360> wl<359> wl<358> wl<357> wl<356> wl<355> wl<354>
+wl<353> wl<352> wl<351> wl<350> wl<349> wl<348> wl<347> wl<346> wl<345>
+wl<344> wl<343> wl<342> wl<341> wl<340> wl<339> wl<338> wl<337> wl<336>
+wl<335> wl<334> wl<333> wl<332> wl<331> wl<330> wl<329> wl<328> wl<327>
+wl<326> wl<325> wl<324> wl<323> wl<322> wl<321> wl<320> wl<319> wl<318>
+wl<317> wl<316> wl<315> wl<314> wl<313> wl<312> wl<311> wl<310> wl<309>
+wl<308> wl<307> wl<306> wl<305> wl<304> wl<303> wl<302> wl<301> wl<300>
+wl<299> wl<298> wl<297> wl<296> wl<295> wl<294> wl<293> wl<292> wl<291>
+wl<290> wl<289> wl<288> wl<287> wl<286> wl<285> wl<284> wl<283> wl<282>
+wl<281> wl<280> wl<279> wl<278> wl<277> wl<276> wl<275> wl<274> wl<273>
+wl<272> wl<271> wl<270> wl<269> wl<268> wl<267> wl<266> wl<265> wl<264>
+wl<263> wl<262> wl<261> wl<260> wl<259> wl<258> wl<257> wl<256> net108  
+deco7_128
XI64 a<6> a<5> a<4> a<3> a<2> a<1> a<0> net<1> net110 wl<255> wl<254> wl<253>
+wl<252> wl<251> wl<250> wl<249> wl<248> wl<247> wl<246> wl<245> wl<244>
+wl<243> wl<242> wl<241> wl<240> wl<239> wl<238> wl<237> wl<236> wl<235>
+wl<234> wl<233> wl<232> wl<231> wl<230> wl<229> wl<228> wl<227> wl<226>
+wl<225> wl<224> wl<223> wl<222> wl<221> wl<220> wl<219> wl<218> wl<217>
+wl<216> wl<215> wl<214> wl<213> wl<212> wl<211> wl<210> wl<209> wl<208>
+wl<207> wl<206> wl<205> wl<204> wl<203> wl<202> wl<201> wl<200> wl<199>
+wl<198> wl<197> wl<196> wl<195> wl<194> wl<193> wl<192> wl<191> wl<190>
+wl<189> wl<188> wl<187> wl<186> wl<185> wl<184> wl<183> wl<182> wl<181>
+wl<180> wl<179> wl<178> wl<177> wl<176> wl<175> wl<174> wl<173> wl<172>
+wl<171> wl<170> wl<169> wl<168> wl<167> wl<166> wl<165> wl<164> wl<163>
+wl<162> wl<161> wl<160> wl<159> wl<158> wl<157> wl<156> wl<155> wl<154>
+wl<153> wl<152> wl<151> wl<150> wl<149> wl<148> wl<147> wl<146> wl<145>
+wl<144> wl<143> wl<142> wl<141> wl<140> wl<139> wl<138> wl<137> wl<136>
+wl<135> wl<134> wl<133> wl<132> wl<131> wl<130> wl<129> wl<128> net108  
+deco7_128
XI55 pre net112   inv Ln=0.35u Wn=8u M=9 Lp=0.35u Wp=16u
XI54 net112 net110   inv Ln=0.35u Wn=8u M=27 Lp=0.35u Wp=16u
XI79 net106 net108   inv Ln=0.35u Wn=8u M=6 Lp=0.35u Wp=16u
XI80 xvld net106   inv Ln=0.35u Wn=10u M=2 Lp=0.35u Wp=20u
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: delay4
* View Name: schematic
************************************************************************

.SUBCKT delay4 A Y
XI47 net38 net39   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI45 net39 net40   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI44 net40 Y   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI46 A net38   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: rl_sel
* View Name: schematic
************************************************************************

.SUBCKT rl_sel a pre sel xvld
XI41 pre pre_out  inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u

MM14 net28 xvld gnd! vbb! NMOS W=8u L=0.35u M=1
MM13 Y A net28 vbb! NMOS W=8u L=0.35u M=1
MM12 Y A vddh2! vddh2! PMOS W=4u L=0.35u M=1.0
MM11 Y xvld vddh2! vddh2! PMOS W=4u L=0.35u M=1.0

MM15 i1 Y gnd! vbb! NMOS W=14u L=350.00n M=1
MM6  i1 Y vddh2! vddh2! PMOS W=28u L=350.00n M=1.0
MM16 i2 i1 gnd! vbb! NMOS W=14u L=350.00n M=1
MM7  i2 i1 vddh2! vddh2! PMOS W=28u L=350.00n M=1.0
MM17 sel i2 gnd! vbb! NMOS W=14u L=350.00n M=1
MM8  sel i2 vddh2! vddh2! PMOS W=28u L=350.00n M=1.0
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: delay6
* View Name: schematic
************************************************************************

.SUBCKT delay6 A Y
XI47 net38 net39   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI45 net39 net40   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI51 net40 net12   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI52 net9 Y   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI46 A net38   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI50 net12 net9   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: sen_ena
* View Name: schematic
************************************************************************

.SUBCKT sen_ena n_ena p_ena xvald
XI70 xvald net25   delay6
XI81 net35 p_ena   inv Ln=0.35u Wn=10u M=9 Lp=0.35u Wp=20u
XI69 net25 net18   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI82 net29 n_ena   inv Ln=0.35u Wn=10u M=9 Lp=0.35u Wp=20u
XI83 net64 net29   inv Ln=0.35u Wn=10u M=3 Lp=0.35u Wp=20u
XI84 net18 net64   inv Ln=0.35u Wn=10u M=1 Lp=0.35u Wp=20u
XI80 net18 net35   inv Ln=0.35u Wn=10u M=2 Lp=0.35u Wp=20u
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: delay16
* View Name: schematic
************************************************************************

.SUBCKT delay16 A Y
XI60 net20 net24   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI47 net15 net39   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI57 net8 net25   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI61 net24 net22   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI59 net25 net26   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI62 net26 net20   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI58 net22 net28   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI63 net28 Y   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI45 net39 net40   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI44 net40 net6   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI48 net6 net4   inv Ln=2.5u Wn=1u M=1 Lp=2.5u Wp=1u
XI51 net4 net12   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI52 net9 net29   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI53 net29 net8   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI46 A net15   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
XI50 net12 net9   inv Ln=2u Wn=1u M=1 Lp=2u Wp=1u
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: xvald
* View Name: schematic
************************************************************************

.SUBCKT xvald pre xvald
XI82 net65 net27   delay6
XI70 net25 net65   delay16
XI24 net27 net28 net22 net25   nand3 Lp=0.35u Wp=3.5u Ln=0.35u Wn=5u
XI17 net28 net27 net21   nand2 Lp=0.35u Wp=3.5u Ln=0.35u Wn=3.5u
XI19 net25 pre net22   nand2 Lp=0.35u Wp=3.5u Ln=0.35u Wn=3.5u
XI18 net22 net21 net28   nand2 Lp=0.35u Wp=3.5u Ln=0.35u Wn=3.5u
XI69 net25 xvald   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
.ENDS

************************************************************************
* Library Name: Lassen_DRAMB
* Cell Name: ctrl256kbm
* View Name: schematic
************************************************************************

.SUBCKT ctrl256kbm a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8>
+a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> cs<511> cs<510> cs<509> cs<508>
+cs<507> cs<506> cs<505> cs<504> cs<503> cs<502> cs<501> cs<500> cs<499>
+cs<498> cs<497> cs<496> cs<495> cs<494> cs<493> cs<492> cs<491> cs<490>
+cs<489> cs<488> cs<487> cs<486> cs<485> cs<484> cs<483> cs<482> cs<481>
+cs<480> cs<479> cs<478> cs<477> cs<476> cs<475> cs<474> cs<473> cs<472>
+cs<471> cs<470> cs<469> cs<468> cs<467> cs<466> cs<465> cs<464> cs<463>
+cs<462> cs<461> cs<460> cs<459> cs<458> cs<457> cs<456> cs<455> cs<454>
+cs<453> cs<452> cs<451> cs<450> cs<449> cs<448> cs<447> cs<446> cs<445>
+cs<444> cs<443> cs<442> cs<441> cs<440> cs<439> cs<438> cs<437> cs<436>
+cs<435> cs<434> cs<433> cs<432> cs<431> cs<430> cs<429> cs<428> cs<427>
+cs<426> cs<425> cs<424> cs<423> cs<422> cs<421> cs<420> cs<419> cs<418>
+cs<417> cs<416> cs<415> cs<414> cs<413> cs<412> cs<411> cs<410> cs<409>
+cs<408> cs<407> cs<406> cs<405> cs<404> cs<403> cs<402> cs<401> cs<400>
+cs<399> cs<398> cs<397> cs<396> cs<395> cs<394> cs<393> cs<392> cs<391>
+cs<390> cs<389> cs<388> cs<387> cs<386> cs<385> cs<384> cs<383> cs<382>
+cs<381> cs<380> cs<379> cs<378> cs<377> cs<376> cs<375> cs<374> cs<373>
+cs<372> cs<371> cs<370> cs<369> cs<368> cs<367> cs<366> cs<365> cs<364>
+cs<363> cs<362> cs<361> cs<360> cs<359> cs<358> cs<357> cs<356> cs<355>
+cs<354> cs<353> cs<352> cs<351> cs<350> cs<349> cs<348> cs<347> cs<346>
+cs<345> cs<344> cs<343> cs<342> cs<341> cs<340> cs<339> cs<338> cs<337>
+cs<336> cs<335> cs<334> cs<333> cs<332> cs<331> cs<330> cs<329> cs<328>
+cs<327> cs<326> cs<325> cs<324> cs<323> cs<322> cs<321> cs<320> cs<319>
+cs<318> cs<317> cs<316> cs<315> cs<314> cs<313> cs<312> cs<311> cs<310>
+cs<309> cs<308> cs<307> cs<306> cs<305> cs<304> cs<303> cs<302> cs<301>
+cs<300> cs<299> cs<298> cs<297> cs<296> cs<295> cs<294> cs<293> cs<292>
+cs<291> cs<290> cs<289> cs<288> cs<287> cs<286> cs<285> cs<284> cs<283>
+cs<282> cs<281> cs<280> cs<279> cs<278> cs<277> cs<276> cs<275> cs<274>
+cs<273> cs<272> cs<271> cs<270> cs<269> cs<268> cs<267> cs<266> cs<265>
+cs<264> cs<263> cs<262> cs<261> cs<260> cs<259> cs<258> cs<257> cs<256>
+cs<255> cs<254> cs<253> cs<252> cs<251> cs<250> cs<249> cs<248> cs<247>
+cs<246> cs<245> cs<244> cs<243> cs<242> cs<241> cs<240> cs<239> cs<238>
+cs<237> cs<236> cs<235> cs<234> cs<233> cs<232> cs<231> cs<230> cs<229>
+cs<228> cs<227> cs<226> cs<225> cs<224> cs<223> cs<222> cs<221> cs<220>
+cs<219> cs<218> cs<217> cs<216> cs<215> cs<214> cs<213> cs<212> cs<211>
+cs<210> cs<209> cs<208> cs<207> cs<206> cs<205> cs<204> cs<203> cs<202>
+cs<201> cs<200> cs<199> cs<198> cs<197> cs<196> cs<195> cs<194> cs<193>
+cs<192> cs<191> cs<190> cs<189> cs<188> cs<187> cs<186> cs<185> cs<184>
+cs<183> cs<182> cs<181> cs<180> cs<179> cs<178> cs<177> cs<176> cs<175>
+cs<174> cs<173> cs<172> cs<171> cs<170> cs<169> cs<168> cs<167> cs<166>
+cs<165> cs<164> cs<163> cs<162> cs<161> cs<160> cs<159> cs<158> cs<157>
+cs<156> cs<155> cs<154> cs<153> cs<152> cs<151> cs<150> cs<149> cs<148>
+cs<147> cs<146> cs<145> cs<144> cs<143> cs<142> cs<141> cs<140> cs<139>
+cs<138> cs<137> cs<136> cs<135> cs<134> cs<133> cs<132> cs<131> cs<130>
+cs<129> cs<128> cs<127> cs<126> cs<125> cs<124> cs<123> cs<122> cs<121>
+cs<120> cs<119> cs<118> cs<117> cs<116> cs<115> cs<114> cs<113> cs<112>
+cs<111> cs<110> cs<109> cs<108> cs<107> cs<106> cs<105> cs<104> cs<103>
+cs<102> cs<101> cs<100> cs<99> cs<98> cs<97> cs<96> cs<95> cs<94> cs<93>
+cs<92> cs<91> cs<90> cs<89> cs<88> cs<87> cs<86> cs<85> cs<84> cs<83> cs<82>
+cs<81> cs<80> cs<79> cs<78> cs<77> cs<76> cs<75> cs<74> cs<73> cs<72> cs<71>
+cs<70> cs<69> cs<68> cs<67> cs<66> cs<65> cs<64> cs<63> cs<62> cs<61> cs<60>
+cs<59> cs<58> cs<57> cs<56> cs<55> cs<54> cs<53> cs<52> cs<51> cs<50> cs<49>
+cs<48> cs<47> cs<46> cs<45> cs<44> cs<43> cs<42> cs<41> cs<40> cs<39> cs<38>
+cs<37> cs<36> cs<35> cs<34> cs<33> cs<32> cs<31> cs<30> cs<29> cs<28> cs<27>
+cs<26> cs<25> cs<24> cs<23> cs<22> cs<21> cs<20> cs<19> cs<18> cs<17> cs<16>
+cs<15> cs<14> cs<13> cs<12> cs<11> cs<10> cs<9> cs<8> cs<7> cs<6> cs<5> cs<4>
+cs<3> cs<2> cs<1> cs<0> ena l_sel main_ena n_ena p_ena pre r_sel w_ wl<511>
+wl<510> wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502>
+wl<501> wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493>
+wl<492> wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484>
+wl<483> wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475>
+wl<474> wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466>
+wl<465> wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457>
+wl<456> wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448>
+wl<447> wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439>
+wl<438> wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430>
+wl<429> wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421>
+wl<420> wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412>
+wl<411> wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403>
+wl<402> wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394>
+wl<393> wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385>
+wl<384> wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376>
+wl<375> wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367>
+wl<366> wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358>
+wl<357> wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349>
+wl<348> wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340>
+wl<339> wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331>
+wl<330> wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322>
+wl<321> wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313>
+wl<312> wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304>
+wl<303> wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295>
+wl<294> wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286>
+wl<285> wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277>
+wl<276> wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268>
+wl<267> wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259>
+wl<258> wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250>
+wl<249> wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241>
+wl<240> wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232>
+wl<231> wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223>
+wl<222> wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214>
+wl<213> wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205>
+wl<204> wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196>
+wl<195> wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187>
+wl<186> wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178>
+wl<177> wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169>
+wl<168> wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160>
+wl<159> wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151>
+wl<150> wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142>
+wl<141> wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133>
+wl<132> wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124>
+wl<123> wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115>
+wl<114> wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106>
+wl<105> wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96>
+wl<95> wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85>
+wl<84> wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74>
+wl<73> wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63>
+wl<62> wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52>
+wl<51> wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41>
+wl<40> wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30>
+wl<29> wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19>
+wl<18> wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8>
+wl<7> wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>
XI139 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> ena w_ net107   atd18m
XI88 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> cs<511> cs<510>
+cs<509> cs<508> cs<507> cs<506> cs<505> cs<504> cs<503> cs<502> cs<501>
+cs<500> cs<499> cs<498> cs<497> cs<496> cs<495> cs<494> cs<493> cs<492>
+cs<491> cs<490> cs<489> cs<488> cs<487> cs<486> cs<485> cs<484> cs<483>
+cs<482> cs<481> cs<480> cs<479> cs<478> cs<477> cs<476> cs<475> cs<474>
+cs<473> cs<472> cs<471> cs<470> cs<469> cs<468> cs<467> cs<466> cs<465>
+cs<464> cs<463> cs<462> cs<461> cs<460> cs<459> cs<458> cs<457> cs<456>
+cs<455> cs<454> cs<453> cs<452> cs<451> cs<450> cs<449> cs<448> cs<447>
+cs<446> cs<445> cs<444> cs<443> cs<442> cs<441> cs<440> cs<439> cs<438>
+cs<437> cs<436> cs<435> cs<434> cs<433> cs<432> cs<431> cs<430> cs<429>
+cs<428> cs<427> cs<426> cs<425> cs<424> cs<423> cs<422> cs<421> cs<420>
+cs<419> cs<418> cs<417> cs<416> cs<415> cs<414> cs<413> cs<412> cs<411>
+cs<410> cs<409> cs<408> cs<407> cs<406> cs<405> cs<404> cs<403> cs<402>
+cs<401> cs<400> cs<399> cs<398> cs<397> cs<396> cs<395> cs<394> cs<393>
+cs<392> cs<391> cs<390> cs<389> cs<388> cs<387> cs<386> cs<385> cs<384>
+cs<383> cs<382> cs<381> cs<380> cs<379> cs<378> cs<377> cs<376> cs<375>
+cs<374> cs<373> cs<372> cs<371> cs<370> cs<369> cs<368> cs<367> cs<366>
+cs<365> cs<364> cs<363> cs<362> cs<361> cs<360> cs<359> cs<358> cs<357>
+cs<356> cs<355> cs<354> cs<353> cs<352> cs<351> cs<350> cs<349> cs<348>
+cs<347> cs<346> cs<345> cs<344> cs<343> cs<342> cs<341> cs<340> cs<339>
+cs<338> cs<337> cs<336> cs<335> cs<334> cs<333> cs<332> cs<331> cs<330>
+cs<329> cs<328> cs<327> cs<326> cs<325> cs<324> cs<323> cs<322> cs<321>
+cs<320> cs<319> cs<318> cs<317> cs<316> cs<315> cs<314> cs<313> cs<312>
+cs<311> cs<310> cs<309> cs<308> cs<307> cs<306> cs<305> cs<304> cs<303>
+cs<302> cs<301> cs<300> cs<299> cs<298> cs<297> cs<296> cs<295> cs<294>
+cs<293> cs<292> cs<291> cs<290> cs<289> cs<288> cs<287> cs<286> cs<285>
+cs<284> cs<283> cs<282> cs<281> cs<280> cs<279> cs<278> cs<277> cs<276>
+cs<275> cs<274> cs<273> cs<272> cs<271> cs<270> cs<269> cs<268> cs<267>
+cs<266> cs<265> cs<264> cs<263> cs<262> cs<261> cs<260> cs<259> cs<258>
+cs<257> cs<256> cs<255> cs<254> cs<253> cs<252> cs<251> cs<250> cs<249>
+cs<248> cs<247> cs<246> cs<245> cs<244> cs<243> cs<242> cs<241> cs<240>
+cs<239> cs<238> cs<237> cs<236> cs<235> cs<234> cs<233> cs<232> cs<231>
+cs<230> cs<229> cs<228> cs<227> cs<226> cs<225> cs<224> cs<223> cs<222>
+cs<221> cs<220> cs<219> cs<218> cs<217> cs<216> cs<215> cs<214> cs<213>
+cs<212> cs<211> cs<210> cs<209> cs<208> cs<207> cs<206> cs<205> cs<204>
+cs<203> cs<202> cs<201> cs<200> cs<199> cs<198> cs<197> cs<196> cs<195>
+cs<194> cs<193> cs<192> cs<191> cs<190> cs<189> cs<188> cs<187> cs<186>
+cs<185> cs<184> cs<183> cs<182> cs<181> cs<180> cs<179> cs<178> cs<177>
+cs<176> cs<175> cs<174> cs<173> cs<172> cs<171> cs<170> cs<169> cs<168>
+cs<167> cs<166> cs<165> cs<164> cs<163> cs<162> cs<161> cs<160> cs<159>
+cs<158> cs<157> cs<156> cs<155> cs<154> cs<153> cs<152> cs<151> cs<150>
+cs<149> cs<148> cs<147> cs<146> cs<145> cs<144> cs<143> cs<142> cs<141>
+cs<140> cs<139> cs<138> cs<137> cs<136> cs<135> cs<134> cs<133> cs<132>
+cs<131> cs<130> cs<129> cs<128> cs<127> cs<126> cs<125> cs<124> cs<123>
+cs<122> cs<121> cs<120> cs<119> cs<118> cs<117> cs<116> cs<115> cs<114>
+cs<113> cs<112> cs<111> cs<110> cs<109> cs<108> cs<107> cs<106> cs<105>
+cs<104> cs<103> cs<102> cs<101> cs<100> cs<99> cs<98> cs<97> cs<96> cs<95>
+cs<94> cs<93> cs<92> cs<91> cs<90> cs<89> cs<88> cs<87> cs<86> cs<85> cs<84>
+cs<83> cs<82> cs<81> cs<80> cs<79> cs<78> cs<77> cs<76> cs<75> cs<74> cs<73>
+cs<72> cs<71> cs<70> cs<69> cs<68> cs<67> cs<66> cs<65> cs<64> cs<63> cs<62>
+cs<61> cs<60> cs<59> cs<58> cs<57> cs<56> cs<55> cs<54> cs<53> cs<52> cs<51>
+cs<50> cs<49> cs<48> cs<47> cs<46> cs<45> cs<44> cs<43> cs<42> cs<41> cs<40>
+cs<39> cs<38> cs<37> cs<36> cs<35> cs<34> cs<33> cs<32> cs<31> cs<30> cs<29>
+cs<28> cs<27> cs<26> cs<25> cs<24> cs<23> cs<22> cs<21> cs<20> cs<19> cs<18>
+cs<17> cs<16> cs<15> cs<14> cs<13> cs<12> cs<11> cs<10> cs<9> cs<8> cs<7>
+cs<6> cs<5> cs<4> cs<3> cs<2> cs<1> cs<0> ena pre net102   col_sel9_512
XI58 a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> ena net107 wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0> xvld   deco9_512
XI99 net102 net75   delay4
XI97 xvld net77 net106 w_   ctg Lp=0.35u Wp=1.4u Ln=0.35u Wn=1.4u
XI96 net85 net77 w_ net106   ctg Lp=0.35u Wp=1.4u Ln=0.35u Wn=1.4u
XI90 xvld net85   delay10
XI146 net116 pre r_sel xvld   rl_sel
XI145 a<8> pre l_sel xvld   rl_sel
XI82 n_ena p_ena xvld   sen_ena
XI100 net75 net98   inv Ln=0.35u Wn=3.5u M=1 Lp=0.35u Wp=7u
XI101 net98 main_ena   inv Ln=0.35u Wn=3.5u M=3 Lp=0.35u Wp=7u
XI95 net104 net102   inv Ln=0.35u Wn=3.5u M=3 Lp=0.35u Wp=7u
XI94 net77 net104   inv Ln=0.35u Wn=3.5u M=1 Lp=0.35u Wp=7u
XI98 w_ net106   inv Ln=0.35u Wn=3.5u M=1 Lp=0.35u Wp=7u
XI108 net107 net108   inv Ln=0.35u Wn=36u M=2 Lp=0.35u Wp=72u
XI81 net114 xvld   inv Ln=0.35u Wn=10u M=9 Lp=0.35u Wp=20u
XI110 net108 pre   inv Ln=0.35u Wn=36u M=5 Lp=0.35u Wp=72u
XI80 net113 net114   inv Ln=0.35u Wn=10u M=3 Lp=0.35u Wp=20u
XI147 a<8> net116   inv Ln=0.35u Wn=3.5u M=1 Lp=0.35u Wp=7u
XI79 pre net113   xvald
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: mc
* View Name: schematic
************************************************************************

.SUBCKT mc bl hv wl
MM0 bl wl cs vbb! NMOS W=700.0n L=350.00n M=1
CC1 cs hv 50f $[CP]
.ENDS

************************************************************************
* Library Name: Lassen_DRAMB
* Cell Name: sa_pre
* View Name: schematic
************************************************************************

.SUBCKT sa_pre bl blb br brb cs io io_ l_sel n_ena p_ena pre r_sel
MM11 net51 net40 net039 vdd! PMOS W=14u L=350.00n M=1
MM15 net40 net51 net039 vdd! PMOS W=14u L=350.00n M=1
MM12 vdd! p_ena net039 vdd! PMOS W=14u L=350.00n M=1
MM80 bl pre blb vbb! NMOS W=1.4u L=350.00n M=1
MM81 vddh! pre blb vbb! NMOS W=1.4u L=350.00n M=1
MM82 vddh! pre bl vbb! NMOS W=1.4u L=350.00n M=1
MM73 br pre brb vbb! NMOS W=1.4u L=350.00n M=1
MM72 vddh! pre br vbb! NMOS W=1.4u L=350.00n M=1
MM71 vddh! pre brb vbb! NMOS W=1.4u L=350.00n M=1
MM76 net40 pre net51 vbb! NMOS W=1.4u L=350.00n M=1
MM75 vddh! pre net40 vbb! NMOS W=1.4u L=350.00n M=1
MM0 blb l_sel net51 vbb! NMOS W=1.4u L=350.00n M=1
MM1 bl l_sel net40 vbb! NMOS W=1.4u L=350.00n M=1
MM77 net51 net40 net081 vbb! NMOS W=7u L=350.00n M=1
MM78 net081 n_ena gnd! vbb! NMOS W=7u L=350.00n M=1
MM79 net40 net51 net081 vbb! NMOS W=7u L=350.00n M=1
MM7 net40 r_sel br vbb! NMOS W=1.4u L=350.00n M=1
MM8 net51 r_sel brb vbb! NMOS W=1.4u L=350.00n M=1
MM9 net40 cs io vbb! NMOS W=1.4u L=350.00n M=1
MM10 io_ cs net51 vbb! NMOS W=1.4u L=350.00n M=1
MM74 vddh! pre net51 vbb! NMOS W=1.4u L=350.00n M=1
.ENDS

************************************************************************
* Library Name: Lassen_DRAMB
* Cell Name: array512x1
* View Name: schematic
************************************************************************

.SUBCKT array512x1 cs io io_ l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>
XI817 bl vddh! wl<307>   mc
XI584 br vddh! wl<133>   mc
XI607 blb vddh! wl<388>   mc
XI813 bl vddh! wl<309>   mc
XI585 brb vddh! wl<128>   mc
XI662 blb vddh! wl<490>   mc
XI680 blb vddh! wl<508>   mc
XI579 br vddh! wl<129>   mc
XI636 bl vddh! wl<447>   mc
XI586 brb vddh! wl<130>   mc
XI639 blb vddh! wl<442>   mc
XI653 blb vddh! wl<428>   mc
XI763 bl vddh! wl<381>   mc
XI587 br vddh! wl<141>   mc
XI757 blb vddh! wl<374>   mc
XI488 brb vddh! wl<220>   mc
XI511 brb vddh! wl<250>   mc
XI582 brb vddh! wl<132>   mc
XI828 bl vddh! wl<287>   mc
XI519 br vddh! wl<231>   mc
XI588 br vddh! wl<143>   mc
XI741 bl vddh! wl<345>   mc
XI789 bl vddh! wl<297>   mc
XI559 brb vddh! wl<180>   mc
XI577 brb vddh! wl<152>   mc
XI578 br vddh! wl<155>   mc
XI567 br vddh! wl<151>   mc
XI589 brb vddh! wl<140>   mc
XI645 blb vddh! wl<422>   mc
XI838 blb vddh! wl<260>   mc
XI661 bl vddh! wl<489>   mc
XI580 br vddh! wl<131>   mc
XI850 bl vddh! wl<267>   mc
XI576 br vddh! wl<153>   mc
XI581 brb vddh! wl<134>   mc
XI583 br vddh! wl<135>   mc
XI575 brb vddh! wl<154>   mc
XI613 bl vddh! wl<409>   mc
XI748 blb vddh! wl<336>   mc
XI535 brb vddh! wl<174>   mc
XI753 bl vddh! wl<339>   mc
XI772 bl vddh! wl<355>   mc
XI833 blb vddh! wl<280>   mc
XI562 br vddh! wl<177>   mc
XI660 blb vddh! wl<488>   mc
XI570 brb vddh! wl<146>   mc
XI538 br vddh! wl<173>   mc
XI548 brb vddh! wl<184>   mc
XI529 brb vddh! wl<232>   mc
XI708 bl vddh! wl<451>   mc
XI668 blb vddh! wl<480>   mc
XI733 bl vddh! wl<325>   mc
XI756 bl vddh! wl<371>   mc
XI549 br vddh! wl<185>   mc
XI805 bl vddh! wl<313>   mc
XI551 brb vddh! wl<190>   mc
XI779 bl vddh! wl<365>   mc
XI539 brb vddh! wl<162>   mc
XI550 brb vddh! wl<186>   mc
XI530 br vddh! wl<235>   mc
XI563 br vddh! wl<145>   mc
XI612 blb vddh! wl<408>   mc
XI571 br vddh! wl<157>   mc
XI724 blb vddh! wl<328>   mc
XI652 bl vddh! wl<431>   mc
XI717 blb vddh! wl<460>   mc
XI764 bl vddh! wl<383>   mc
XI545 br vddh! wl<163>   mc
XI787 bl vddh! wl<299>   mc
XI536 brb vddh! wl<172>   mc
XI544 brb vddh! wl<166>   mc
XI527 brb vddh! wl<234>   mc
XI684 blb vddh! wl<496>   mc
XI693 blb vddh! wl<470>   mc
XI561 br vddh! wl<179>   mc
XI644 bl vddh! wl<419>   mc
XI569 brb vddh! wl<144>   mc
XI537 br vddh! wl<175>   mc
XI546 br vddh! wl<161>   mc
XI528 br vddh! wl<233>   mc
XI740 blb vddh! wl<344>   mc
XI547 br vddh! wl<187>   mc
XI796 blb vddh! wl<288>   mc
XI560 brb vddh! wl<182>   mc
XI568 br vddh! wl<149>   mc
XI700 bl vddh! wl<479>   mc
XI827 bl vddh! wl<285>   mc
XI677 bl vddh! wl<505>   mc
XI566 brb vddh! wl<148>   mc
XI557 br vddh! wl<181>   mc
XI629 blb vddh! wl<438>   mc
XI542 br vddh! wl<167>   mc
XI716 bl vddh! wl<463>   mc
XI533 br vddh! wl<169>   mc
XI685 bl vddh! wl<501>   mc
XI556 brb vddh! wl<176>   mc
XI573 brb vddh! wl<156>   mc
XI816 blb vddh! wl<310>   mc
XI732 blb vddh! wl<320>   mc
XI798 bl vddh! wl<295>   mc
XI849 blb vddh! wl<264>   mc
XI676 blb vddh! wl<504>   mc
XI543 brb vddh! wl<164>   mc
XI692 bl vddh! wl<467>   mc
XI534 brb vddh! wl<170>   mc
XI701 blb vddh! wl<476>   mc
XI558 br vddh! wl<183>   mc
XI574 brb vddh! wl<158>   mc
XI553 br vddh! wl<191>   mc
XI781 blb vddh! wl<364>   mc
XI540 brb vddh! wl<160>   mc
XI552 brb vddh! wl<188>   mc
XI531 br vddh! wl<171>   mc
XI709 blb vddh! wl<454>   mc
XI554 br vddh! wl<189>   mc
XI605 bl vddh! wl<389>   mc
XI565 brb vddh! wl<150>   mc
XI555 brb vddh! wl<178>   mc
XI541 br vddh! wl<165>   mc
XI532 brb vddh! wl<168>   mc
XI837 blb vddh! wl<262>   mc
XI620 blb vddh! wl<400>   mc
XI807 blb vddh! wl<318>   mc
XI564 br vddh! wl<147>   mc
XI604 blb vddh! wl<384>   mc
XI572 br vddh! wl<159>   mc
XI725 bl vddh! wl<329>   mc
XI628 bl vddh! wl<435>   mc
XI621 bl vddh! wl<405>   mc
XI690 bl vddh! wl<497>   mc
XI754 bl vddh! wl<337>   mc
XI516 br vddh! wl<227>   mc
XI730 bl vddh! wl<333>   mc
XI524 br vddh! wl<239>   mc
XI691 bl vddh! wl<465>   mc
XI507 br vddh! wl<253>   mc
XI486 brb vddh! wl<218>   mc
XI493 br vddh! wl<213>   mc
XI506 brb vddh! wl<242>   mc
XI659 bl vddh! wl<491>   mc
XI517 brb vddh! wl<230>   mc
XI618 bl vddh! wl<413>   mc
XI525 brb vddh! wl<236>   mc
XI714 blb vddh! wl<450>   mc
XI738 bl vddh! wl<321>   mc
XI492 brb vddh! wl<208>   mc
XI504 br vddh! wl<245>   mc
XI667 blb vddh! wl<482>   mc
XI731 blb vddh! wl<322>   mc
XI505 brb vddh! wl<240>   mc
XI485 br vddh! wl<217>   mc
XI847 blb vddh! wl<266>   mc
XI510 brb vddh! wl<254>   mc
XI746 bl vddh! wl<349>   mc
XI495 brb vddh! wl<212>   mc
XI626 bl vddh! wl<401>   mc
XI611 bl vddh! wl<411>   mc
XI699 bl vddh! wl<477>   mc
XI610 bl vddh! wl<385>   mc
XI675 bl vddh! wl<507>   mc
XI487 brb vddh! wl<222>   mc
XI825 blb vddh! wl<272>   mc
XI602 bl vddh! wl<397>   mc
XI762 blb vddh! wl<370>   mc
XI494 br vddh! wl<215>   mc
XI508 br vddh! wl<255>   mc
XI651 bl vddh! wl<429>   mc
XI518 brb vddh! wl<228>   mc
XI509 brb vddh! wl<252>   mc
XI526 brb vddh! wl<238>   mc
XI650 blb vddh! wl<418>   mc
XI683 blb vddh! wl<498>   mc
XI814 bl vddh! wl<311>   mc
XI512 br vddh! wl<249>   mc
XI707 bl vddh! wl<449>   mc
XI520 br vddh! wl<229>   mc
XI499 br vddh! wl<241>   mc
XI482 br vddh! wl<193>   mc
XI603 blb vddh! wl<386>   mc
XI498 br vddh! wl<209>   mc
XI513 brb vddh! wl<248>   mc
XI722 bl vddh! wl<459>   mc
XI521 brb vddh! wl<224>   mc
XI658 bl vddh! wl<427>   mc
XI723 bl vddh! wl<331>   mc
XI835 bl vddh! wl<257>   mc
XI627 bl vddh! wl<433>   mc
XI496 brb vddh! wl<214>   mc
XI826 blb vddh! wl<274>   mc
XI489 br vddh! wl<223>   mc
XI497 br vddh! wl<211>   mc
XI481 br vddh! wl<195>   mc
XI642 bl vddh! wl<443>   mc
XI698 blb vddh! wl<466>   mc
XI515 br vddh! wl<225>   mc
XI674 bl vddh! wl<481>   mc
XI523 br vddh! wl<237>   mc
XI491 brb vddh! wl<210>   mc
XI502 brb vddh! wl<244>   mc
XI643 bl vddh! wl<417>   mc
XI715 bl vddh! wl<461>   mc
XI503 br vddh! wl<247>   mc
XI484 brb vddh! wl<216>   mc
XI619 blb vddh! wl<402>   mc
XI501 brb vddh! wl<246>   mc
XI483 br vddh! wl<219>   mc
XI666 bl vddh! wl<493>   mc
XI706 bl vddh! wl<475>   mc
XI490 br vddh! wl<221>   mc
XI500 br vddh! wl<243>   mc
XI514 br vddh! wl<251>   mc
XI682 bl vddh! wl<509>   mc
XI522 brb vddh! wl<226>   mc
XI713 blb vddh! wl<448>   mc
XI770 bl vddh! wl<379>   mc
XI702 blb vddh! wl<478>   mc
XI729 bl vddh! wl<335>   mc
XI744 blb vddh! wl<348>   mc
XI649 blb vddh! wl<416>   mc
XI829 blb vddh! wl<284>   mc
XI760 bl vddh! wl<373>   mc
XI678 blb vddh! wl<506>   mc
XI818 bl vddh! wl<305>   mc
XI820 bl vddh! wl<275>   mc
XI734 bl vddh! wl<327>   mc
XI694 blb vddh! wl<468>   mc
XI705 blb vddh! wl<472>   mc
XI832 bl vddh! wl<281>   mc
XI689 bl vddh! wl<499>   mc
XI841 blb vddh! wl<256>   mc
XI670 bl vddh! wl<487>   mc
XI783 blb vddh! wl<362>   mc
XI726 blb vddh! wl<330>   mc
XI840 bl vddh! wl<261>   mc
XI822 blb vddh! wl<276>   mc
XI615 blb vddh! wl<414>   mc
XI679 blb vddh! wl<510>   mc
XI669 bl vddh! wl<485>   mc
XI804 blb vddh! wl<312>   mc
XI632 bl vddh! wl<437>   mc
XI703 blb vddh! wl<474>   mc
XI322 br vddh! wl<1>   mc
XI371 br vddh! wl<49>   mc
XI819 bl vddh! wl<273>   mc
XI321 br vddh! wl<3>   mc
XI782 blb vddh! wl<366>   mc
XI594 br vddh! wl<139>   mc
XI808 blb vddh! wl<316>   mc
XI593 brb vddh! wl<136>   mc
XI799 blb vddh! wl<292>   mc
XI592 br vddh! wl<137>   mc
XI790 blb vddh! wl<298>   mc
XI591 brb vddh! wl<138>   mc
XI749 bl vddh! wl<341>   mc
XI590 brb vddh! wl<142>   mc
XI765 blb vddh! wl<380>   mc
XI403 br vddh! wl<107>   mc
XI405 br vddh! wl<105>   mc
XI406 brb vddh! wl<106>   mc
XI407 brb vddh! wl<110>   mc
XI408 brb vddh! wl<108>   mc
XI409 br vddh! wl<111>   mc
XI411 brb vddh! wl<98>   mc
XI410 br vddh! wl<109>   mc
XI412 brb vddh! wl<96>   mc
XI413 br vddh! wl<101>   mc
XI414 br vddh! wl<103>   mc
XI415 brb vddh! wl<100>   mc
XI416 brb vddh! wl<102>   mc
XI417 br vddh! wl<99>   mc
XI418 br vddh! wl<97>   mc
XI420 brb vddh! wl<120>   mc
XI419 br vddh! wl<123>   mc
XI422 brb vddh! wl<122>   mc
XI421 br vddh! wl<121>   mc
XI423 brb vddh! wl<126>   mc
XI424 brb vddh! wl<124>   mc
XI425 br vddh! wl<127>   mc
XI426 br vddh! wl<125>   mc
XI427 brb vddh! wl<114>   mc
XI428 brb vddh! wl<112>   mc
XI429 br vddh! wl<117>   mc
XI430 br vddh! wl<119>   mc
XI402 br vddh! wl<43>   mc
XI401 brb vddh! wl<40>   mc
XI400 br vddh! wl<41>   mc
XI399 brb vddh! wl<42>   mc
XI398 brb vddh! wl<46>   mc
XI397 brb vddh! wl<44>   mc
XI310 brb vddh! wl<10>   mc
XI431 brb vddh! wl<116>   mc
XI396 br vddh! wl<47>   mc
XI801 bl vddh! wl<291>   mc
XI784 bl vddh! wl<361>   mc
XI395 br vddh! wl<45>   mc
XI735 blb vddh! wl<324>   mc
XI768 bl vddh! wl<377>   mc
XI663 blb vddh! wl<494>   mc
XI695 bl vddh! wl<471>   mc
XI759 bl vddh! wl<375>   mc
XI317 br vddh! wl<5>   mc
XI319 brb vddh! wl<4>   mc
XI600 blb vddh! wl<396>   mc
XI601 bl vddh! wl<399>   mc
XI655 blb vddh! wl<426>   mc
XI846 blb vddh! wl<270>   mc
XI751 blb vddh! wl<340>   mc
XI834 bl vddh! wl<283>   mc
XI743 blb vddh! wl<350>   mc
XI719 blb vddh! wl<458>   mc
XI792 blb vddh! wl<300>   mc
XI671 blb vddh! wl<484>   mc
XI623 blb vddh! wl<404>   mc
XI810 bl vddh! wl<317>   mc
XI647 bl vddh! wl<423>   mc
XI780 bl vddh! wl<367>   mc
XI475 brb vddh! wl<194>   mc
XI635 bl vddh! wl<445>   mc
XI467 br vddh! wl<203>   mc
XI771 bl vddh! wl<353>   mc
XI769 blb vddh! wl<376>   mc
XI806 blb vddh! wl<314>   mc
XI476 brb vddh! wl<192>   mc
XI633 blb vddh! wl<432>   mc
XI394 brb vddh! wl<34>   mc
XI393 brb vddh! wl<32>   mc
XI468 brb vddh! wl<200>   mc
XI803 bl vddh! wl<315>   mc
XI794 bl vddh! wl<301>   mc
XI392 br vddh! wl<37>   mc
XI391 br vddh! wl<39>   mc
XI474 br vddh! wl<205>   mc
XI390 brb vddh! wl<36>   mc
XI774 blb vddh! wl<356>   mc
XI755 bl vddh! wl<369>   mc
XI307 br vddh! wl<11>   mc
XI824 bl vddh! wl<277>   mc
XI389 brb vddh! wl<38>   mc
XI795 blb vddh! wl<290>   mc
XI812 blb vddh! wl<304>   mc
XI388 br vddh! wl<35>   mc
XI320 brb vddh! wl<6>   mc
XI387 br vddh! wl<33>   mc
XI598 blb vddh! wl<394>   mc
XI386 br vddh! wl<59>   mc
XI385 brb vddh! wl<56>   mc
XI384 br vddh! wl<57>   mc
XI383 brb vddh! wl<58>   mc
XI381 brb vddh! wl<60>   mc
XI382 brb vddh! wl<62>   mc
XI380 br vddh! wl<63>   mc
XI379 br vddh! wl<61>   mc
XI378 brb vddh! wl<50>   mc
XI377 brb vddh! wl<48>   mc
XI599 blb vddh! wl<398>   mc
XI376 br vddh! wl<53>   mc
XI375 br vddh! wl<55>   mc
XI773 blb vddh! wl<358>   mc
XI374 brb vddh! wl<52>   mc
XI373 brb vddh! wl<54>   mc
XI372 br vddh! wl<51>   mc
XI711 bl vddh! wl<455>   mc
XI786 bl vddh! wl<363>   mc
XI687 blb vddh! wl<500>   mc
XI830 blb vddh! wl<286>   mc
XI739 bl vddh! wl<347>   mc
XI637 blb vddh! wl<444>   mc
XI432 brb vddh! wl<118>   mc
XI638 blb vddh! wl<446>   mc
XI473 br vddh! wl<207>   mc
XI433 br vddh! wl<115>   mc
XI775 bl vddh! wl<359>   mc
XI848 bl vddh! wl<265>   mc
XI641 blb vddh! wl<440>   mc
XI747 blb vddh! wl<338>   mc
XI479 brb vddh! wl<196>   mc
XI823 bl vddh! wl<279>   mc
XI471 brb vddh! wl<206>   mc
XI778 blb vddh! wl<354>   mc
XI844 bl vddh! wl<271>   mc
XI776 bl vddh! wl<357>   mc
XI313 br vddh! wl<15>   mc
XI777 blb vddh! wl<352>   mc
XI434 br vddh! wl<113>   mc
XI435 br vddh! wl<81>   mc
XI480 brb vddh! wl<198>   mc
XI640 bl vddh! wl<441>   mc
XI472 brb vddh! wl<204>   mc
XI767 blb vddh! wl<378>   mc
XI478 br vddh! wl<199>   mc
XI311 brb vddh! wl<14>   mc
XI309 br vddh! wl<9>   mc
XI843 bl vddh! wl<269>   mc
XI314 br vddh! wl<13>   mc
XI470 brb vddh! wl<202>   mc
XI436 br vddh! wl<83>   mc
XI815 blb vddh! wl<308>   mc
XI323 br vddh! wl<27>   mc
XI437 brb vddh! wl<86>   mc
XI788 blb vddh! wl<296>   mc
XI438 brb vddh! wl<84>   mc
XI439 br vddh! wl<87>   mc
XI440 br vddh! wl<85>   mc
XI441 brb vddh! wl<80>   mc
XI442 brb vddh! wl<82>   mc
XI845 blb vddh! wl<268>   mc
XI836 bl vddh! wl<259>   mc
XI797 bl vddh! wl<293>   mc
XI443 br vddh! wl<93>   mc
XI477 br vddh! wl<197>   mc
XI631 bl vddh! wl<439>   mc
XI469 br vddh! wl<201>   mc
XI681 bl vddh! wl<511>   mc
XI821 blb vddh! wl<278>   mc
XI648 bl vddh! wl<421>   mc
XI697 blb vddh! wl<464>   mc
XI315 brb vddh! wl<2>   mc
XI606 bl vddh! wl<391>   mc
XI656 bl vddh! wl<425>   mc
XI758 blb vddh! wl<372>   mc
XI672 blb vddh! wl<486>   mc
XI444 br vddh! wl<95>   mc
XI445 brb vddh! wl<92>   mc
XI324 brb vddh! wl<24>   mc
XI325 br vddh! wl<25>   mc
XI326 brb vddh! wl<26>   mc
XI446 brb vddh! wl<94>   mc
XI447 brb vddh! wl<90>   mc
XI327 brb vddh! wl<30>   mc
XI448 br vddh! wl<89>   mc
XI328 brb vddh! wl<28>   mc
XI616 blb vddh! wl<412>   mc
XI329 br vddh! wl<31>   mc
XI449 brb vddh! wl<88>   mc
XI450 br vddh! wl<91>   mc
XI451 br vddh! wl<65>   mc
XI452 br vddh! wl<67>   mc
XI453 brb vddh! wl<70>   mc
XI454 brb vddh! wl<68>   mc
XI721 blb vddh! wl<456>   mc
XI842 blb vddh! wl<258>   mc
XI664 blb vddh! wl<492>   mc
XI737 bl vddh! wl<323>   mc
XI718 blb vddh! wl<462>   mc
XI831 blb vddh! wl<282>   mc
XI839 bl vddh! wl<263>   mc
XI622 bl vddh! wl<407>   mc
XI455 br vddh! wl<71>   mc
XI745 bl vddh! wl<351>   mc
XI736 blb vddh! wl<326>   mc
XI609 bl vddh! wl<387>   mc
XI330 br vddh! wl<29>   mc
XI331 brb vddh! wl<18>   mc
XI404 brb vddh! wl<104>   mc
XI316 brb vddh! wl<0>   mc
XI654 blb vddh! wl<430>   mc
XI720 bl vddh! wl<457>   mc
XI750 bl vddh! wl<343>   mc
XI696 bl vddh! wl<469>   mc
XI332 brb vddh! wl<16>   mc
XI791 blb vddh! wl<302>   mc
XI614 blb vddh! wl<410>   mc
XI595 bl vddh! wl<395>   mc
XI608 blb vddh! wl<390>   mc
XI333 br vddh! wl<21>   mc
XI308 brb vddh! wl<8>   mc
XI766 blb vddh! wl<382>   mc
XI456 br vddh! wl<69>   mc
XI625 bl vddh! wl<403>   mc
XI596 blb vddh! wl<392>   mc
XI597 bl vddh! wl<393>   mc
XI630 blb vddh! wl<436>   mc
XI634 blb vddh! wl<434>   mc
XI457 brb vddh! wl<64>   mc
XI742 blb vddh! wl<346>   mc
XI761 blb vddh! wl<368>   mc
XI318 br vddh! wl<7>   mc
XI624 blb vddh! wl<406>   mc
XI617 bl vddh! wl<415>   mc
XI809 bl vddh! wl<319>   mc
XI458 brb vddh! wl<66>   mc
XI459 br vddh! wl<77>   mc
XI460 br vddh! wl<79>   mc
XI334 br vddh! wl<23>   mc
XI704 bl vddh! wl<473>   mc
XI657 blb vddh! wl<424>   mc
XI785 blb vddh! wl<360>   mc
XI335 brb vddh! wl<20>   mc
XI461 brb vddh! wl<76>   mc
XI688 blb vddh! wl<502>   mc
XI336 brb vddh! wl<22>   mc
XI337 br vddh! wl<19>   mc
XI686 bl vddh! wl<503>   mc
XI793 bl vddh! wl<303>   mc
XI462 brb vddh! wl<78>   mc
XI338 br vddh! wl<17>   mc
XI710 blb vddh! wl<452>   mc
XI463 brb vddh! wl<74>   mc
XI811 blb vddh! wl<306>   mc
XI646 blb vddh! wl<420>   mc
XI673 bl vddh! wl<483>   mc
XI752 blb vddh! wl<342>   mc
XI728 blb vddh! wl<332>   mc
XI464 br vddh! wl<73>   mc
XI665 bl vddh! wl<495>   mc
XI802 bl vddh! wl<289>   mc
XI712 bl vddh! wl<453>   mc
XI312 brb vddh! wl<12>   mc
XI465 brb vddh! wl<72>   mc
XI466 br vddh! wl<75>   mc
XI727 blb vddh! wl<334>   mc
XI800 blb vddh! wl<294>   mc
XI304 bl blb br brb cs io io_ l_sel n_ena p_ena pre r_sel   sa_pre
CC51 blb gnd! 250f $[CP]
CC52 bl gnd! 250f $[CP]
CC8 brb gnd! 250f $[CP]
CC7 br gnd! 250f $[CP]
.ENDS

************************************************************************
* Library Name: Lassen_DRAMB
* Cell Name: block512x512n
* View Name: schematic
************************************************************************

.SUBCKT block512x512n a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9>
+a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> ena i_o w_
XI102 net696 i_o ena net690   ctg Lp=0.35u Wp=1.4u Ln=0.35u Wn=1.4u
XI100 ena net690   inv Ln=0.35u Wn=1.4u M=1 Lp=0.35u Wp=1.4u
XI1367 a<0> net696 net9403 net9404 main_ena pre w_   io
XI1366 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6>
+a<5> a<4> a<3> a<2> a<1> a<0> cl<511> cl<510> cl<509> cl<508> cl<507> cl<506>
+cl<505> cl<504> cl<503> cl<502> cl<501> cl<500> cl<499> cl<498> cl<497>
+cl<496> cl<495> cl<494> cl<493> cl<492> cl<491> cl<490> cl<489> cl<488>
+cl<487> cl<486> cl<485> cl<484> cl<483> cl<482> cl<481> cl<480> cl<479>
+cl<478> cl<477> cl<476> cl<475> cl<474> cl<473> cl<472> cl<471> cl<470>
+cl<469> cl<468> cl<467> cl<466> cl<465> cl<464> cl<463> cl<462> cl<461>
+cl<460> cl<459> cl<458> cl<457> cl<456> cl<455> cl<454> cl<453> cl<452>
+cl<451> cl<450> cl<449> cl<448> cl<447> cl<446> cl<445> cl<444> cl<443>
+cl<442> cl<441> cl<440> cl<439> cl<438> cl<437> cl<436> cl<435> cl<434>
+cl<433> cl<432> cl<431> cl<430> cl<429> cl<428> cl<427> cl<426> cl<425>
+cl<424> cl<423> cl<422> cl<421> cl<420> cl<419> cl<418> cl<417> cl<416>
+cl<415> cl<414> cl<413> cl<412> cl<411> cl<410> cl<409> cl<408> cl<407>
+cl<406> cl<405> cl<404> cl<403> cl<402> cl<401> cl<400> cl<399> cl<398>
+cl<397> cl<396> cl<395> cl<394> cl<393> cl<392> cl<391> cl<390> cl<389>
+cl<388> cl<387> cl<386> cl<385> cl<384> cl<383> cl<382> cl<381> cl<380>
+cl<379> cl<378> cl<377> cl<376> cl<375> cl<374> cl<373> cl<372> cl<371>
+cl<370> cl<369> cl<368> cl<367> cl<366> cl<365> cl<364> cl<363> cl<362>
+cl<361> cl<360> cl<359> cl<358> cl<357> cl<356> cl<355> cl<354> cl<353>
+cl<352> cl<351> cl<350> cl<349> cl<348> cl<347> cl<346> cl<345> cl<344>
+cl<343> cl<342> cl<341> cl<340> cl<339> cl<338> cl<337> cl<336> cl<335>
+cl<334> cl<333> cl<332> cl<331> cl<330> cl<329> cl<328> cl<327> cl<326>
+cl<325> cl<324> cl<323> cl<322> cl<321> cl<320> cl<319> cl<318> cl<317>
+cl<316> cl<315> cl<314> cl<313> cl<312> cl<311> cl<310> cl<309> cl<308>
+cl<307> cl<306> cl<305> cl<304> cl<303> cl<302> cl<301> cl<300> cl<299>
+cl<298> cl<297> cl<296> cl<295> cl<294> cl<293> cl<292> cl<291> cl<290>
+cl<289> cl<288> cl<287> cl<286> cl<285> cl<284> cl<283> cl<282> cl<281>
+cl<280> cl<279> cl<278> cl<277> cl<276> cl<275> cl<274> cl<273> cl<272>
+cl<271> cl<270> cl<269> cl<268> cl<267> cl<266> cl<265> cl<264> cl<263>
+cl<262> cl<261> cl<260> cl<259> cl<258> cl<257> cl<256> cl<255> cl<254>
+cl<253> cl<252> cl<251> cl<250> cl<249> cl<248> cl<247> cl<246> cl<245>
+cl<244> cl<243> cl<242> cl<241> cl<240> cl<239> cl<238> cl<237> cl<236>
+cl<235> cl<234> cl<233> cl<232> cl<231> cl<230> cl<229> cl<228> cl<227>
+cl<226> cl<225> cl<224> cl<223> cl<222> cl<221> cl<220> cl<219> cl<218>
+cl<217> cl<216> cl<215> cl<214> cl<213> cl<212> cl<211> cl<210> cl<209>
+cl<208> cl<207> cl<206> cl<205> cl<204> cl<203> cl<202> cl<201> cl<200>
+cl<199> cl<198> cl<197> cl<196> cl<195> cl<194> cl<193> cl<192> cl<191>
+cl<190> cl<189> cl<188> cl<187> cl<186> cl<185> cl<184> cl<183> cl<182>
+cl<181> cl<180> cl<179> cl<178> cl<177> cl<176> cl<175> cl<174> cl<173>
+cl<172> cl<171> cl<170> cl<169> cl<168> cl<167> cl<166> cl<165> cl<164>
+cl<163> cl<162> cl<161> cl<160> cl<159> cl<158> cl<157> cl<156> cl<155>
+cl<154> cl<153> cl<152> cl<151> cl<150> cl<149> cl<148> cl<147> cl<146>
+cl<145> cl<144> cl<143> cl<142> cl<141> cl<140> cl<139> cl<138> cl<137>
+cl<136> cl<135> cl<134> cl<133> cl<132> cl<131> cl<130> cl<129> cl<128>
+cl<127> cl<126> cl<125> cl<124> cl<123> cl<122> cl<121> cl<120> cl<119>
+cl<118> cl<117> cl<116> cl<115> cl<114> cl<113> cl<112> cl<111> cl<110>
+cl<109> cl<108> cl<107> cl<106> cl<105> cl<104> cl<103> cl<102> cl<101>
+cl<100> cl<99> cl<98> cl<97> cl<96> cl<95> cl<94> cl<93> cl<92> cl<91> cl<90>
+cl<89> cl<88> cl<87> cl<86> cl<85> cl<84> cl<83> cl<82> cl<81> cl<80> cl<79>
+cl<78> cl<77> cl<76> cl<75> cl<74> cl<73> cl<72> cl<71> cl<70> cl<69> cl<68>
+cl<67> cl<66> cl<65> cl<64> cl<63> cl<62> cl<61> cl<60> cl<59> cl<58> cl<57>
+cl<56> cl<55> cl<54> cl<53> cl<52> cl<51> cl<50> cl<49> cl<48> cl<47> cl<46>
+cl<45> cl<44> cl<43> cl<42> cl<41> cl<40> cl<39> cl<38> cl<37> cl<36> cl<35>
+cl<34> cl<33> cl<32> cl<31> cl<30> cl<29> cl<28> cl<27> cl<26> cl<25> cl<24>
+cl<23> cl<22> cl<21> cl<20> cl<19> cl<18> cl<17> cl<16> cl<15> cl<14> cl<13>
+cl<12> cl<11> cl<10> cl<9> cl<8> cl<7> cl<6> cl<5> cl<4> cl<3> cl<2> cl<1>
+cl<0> ena l_sel main_ena n_ena p_ena pre r_sel w_ wl<511> wl<510> wl<509>
+wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501> wl<500>
+wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492> wl<491>
+wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483> wl<482>
+wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474> wl<473>
+wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465> wl<464>
+wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456> wl<455>
+wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447> wl<446>
+wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438> wl<437>
+wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429> wl<428>
+wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420> wl<419>
+wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411> wl<410>
+wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402> wl<401>
+wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393> wl<392>
+wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384> wl<383>
+wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375> wl<374>
+wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366> wl<365>
+wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357> wl<356>
+wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348> wl<347>
+wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339> wl<338>
+wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330> wl<329>
+wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321> wl<320>
+wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312> wl<311>
+wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303> wl<302>
+wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294> wl<293>
+wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285> wl<284>
+wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276> wl<275>
+wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267> wl<266>
+wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258> wl<257>
+wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249> wl<248>
+wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240> wl<239>
+wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231> wl<230>
+wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222> wl<221>
+wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213> wl<212>
+wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204> wl<203>
+wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195> wl<194>
+wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186> wl<185>
+wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177> wl<176>
+wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168> wl<167>
+wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159> wl<158>
+wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150> wl<149>
+wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141> wl<140>
+wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132> wl<131>
+wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123> wl<122>
+wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114> wl<113>
+wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105> wl<104>
+wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95> wl<94>
+wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84> wl<83>
+wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73> wl<72>
+wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62> wl<61>
+wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51> wl<50>
+wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40> wl<39>
+wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29> wl<28>
+wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18> wl<17>
+wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7> wl<6>
+wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   ctrl256kbm
XI887 cl<34> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI888 cl<38> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI889 cl<44> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI890 cl<39> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI891 cl<37> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI892 cl<36> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI893 cl<45> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI894 cl<47> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI895 cl<46> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI896 cl<42> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI897 cl<43> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI898 cl<41> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI899 cl<40> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI900 cl<56> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI901 cl<57> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI902 cl<59> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI903 cl<58> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI904 cl<62> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI905 cl<63> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI906 cl<61> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI907 cl<60> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI908 cl<52> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI909 cl<53> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI910 cl<55> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI911 cl<54> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI912 cl<50> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI913 cl<51> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI914 cl<49> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI915 cl<48> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI916 cl<32> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI917 cl<33> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI918 cl<97> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI919 cl<96> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI920 cl<112> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI922 cl<115> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI923 cl<114> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI921 cl<113> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI924 cl<118> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI925 cl<119> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI926 cl<117> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI927 cl<116> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI928 cl<124> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI929 cl<125> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI930 cl<127> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI931 cl<126> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI932 cl<122> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI933 cl<123> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI934 cl<121> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI935 cl<120> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI936 cl<104> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI937 cl<105> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI938 cl<107> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI939 cl<106> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI940 cl<110> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI941 cl<111> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI942 cl<109> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI943 cl<100> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI944 cl<101> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI945 cl<103> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI946 cl<108> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI947 cl<102> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI948 cl<98> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI949 cl<99> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI950 cl<67> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI951 cl<66> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI952 cl<70> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI953 cl<76> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI954 cl<71> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI955 cl<69> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI956 cl<68> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI957 cl<77> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI958 cl<79> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI959 cl<78> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI960 cl<74> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI961 cl<75> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI962 cl<73> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI963 cl<72> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI964 cl<88> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI965 cl<89> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI966 cl<91> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI967 cl<90> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI968 cl<94> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI969 cl<95> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI970 cl<93> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI971 cl<92> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI972 cl<84> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI973 cl<85> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI974 cl<87> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI975 cl<86> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI976 cl<82> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI977 cl<83> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI978 cl<81> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI979 cl<80> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI980 cl<64> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI981 cl<65> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI982 cl<193> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI983 cl<192> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI984 cl<208> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI987 cl<210> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI988 cl<214> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI985 cl<209> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI986 cl<211> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI989 cl<215> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI990 cl<213> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI991 cl<212> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI992 cl<220> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI993 cl<221> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI994 cl<223> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI995 cl<222> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI996 cl<219> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI997 cl<218> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI998 cl<217> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI999 cl<216> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1000 cl<200> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1001 cl<201> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1002 cl<203> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1003 cl<202> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1004 cl<206> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1005 cl<207> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1006 cl<205> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1007 cl<196> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1008 cl<197> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1009 cl<199> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1010 cl<204> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1011 cl<198> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1012 cl<194> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1013 cl<195> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1014 cl<227> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1015 cl<226> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1016 cl<230> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1017 cl<236> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1018 cl<231> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1019 cl<229> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1020 cl<228> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1021 cl<237> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1022 cl<239> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1023 cl<238> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1024 cl<234> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1025 cl<235> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1026 cl<233> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1027 cl<232> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1028 cl<248> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1029 cl<249> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1030 cl<251> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1031 cl<250> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1032 cl<254> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1033 cl<255> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1034 cl<253> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1035 cl<252> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1036 cl<244> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1037 cl<245> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1038 cl<247> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1039 cl<246> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1040 cl<242> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1041 cl<243> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1042 cl<241> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1043 cl<240> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1044 cl<224> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1045 cl<225> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1046 cl<161> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1047 cl<160> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1048 cl<176> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1049 cl<177> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1050 cl<179> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1051 cl<178> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1052 cl<182> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1053 cl<183> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1054 cl<181> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1055 cl<180> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1056 cl<188> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1057 cl<189> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1058 cl<191> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1059 cl<190> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1060 cl<186> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1061 cl<187> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1062 cl<185> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1063 cl<184> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1064 cl<168> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1065 cl<169> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1066 cl<171> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1067 cl<170> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1068 cl<174> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1069 cl<175> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1070 cl<173> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1071 cl<164> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1072 cl<165> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1073 cl<167> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1074 cl<172> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1075 cl<166> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1076 cl<162> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1077 cl<163> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1078 cl<131> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1079 cl<130> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1080 cl<134> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1081 cl<140> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1082 cl<135> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1083 cl<133> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1084 cl<132> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1085 cl<141> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1086 cl<143> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1087 cl<142> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1088 cl<138> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1089 cl<139> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1090 cl<137> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1091 cl<136> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1092 cl<152> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1093 cl<153> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1094 cl<155> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1095 cl<154> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1096 cl<158> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1097 cl<159> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1098 cl<157> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1099 cl<156> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1100 cl<148> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1101 cl<149> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1102 cl<151> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1103 cl<150> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1104 cl<146> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1105 cl<147> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1106 cl<145> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1107 cl<144> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1108 cl<128> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1109 cl<129> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1110 cl<385> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1111 cl<384> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1114 cl<403> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI856 cl<3> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI857 cl<2> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI858 cl<6> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI862 cl<12> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI859 cl<7> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI860 cl<5> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI861 cl<4> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI863 cl<13> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI864 cl<15> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI865 cl<14> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI866 cl<10> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI867 cl<11> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI868 cl<9> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI869 cl<8> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI870 cl<24> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI871 cl<25> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI872 cl<27> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI873 cl<26> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI874 cl<30> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI875 cl<31> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI876 cl<29> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI877 cl<28> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI878 cl<20> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI879 cl<21> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI880 cl<23> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI881 cl<22> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI882 cl<18> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI883 cl<19> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI884 cl<17> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI885 cl<16> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1115 cl<402> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1112 cl<400> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1113 cl<401> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1116 cl<406> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1117 cl<407> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1118 cl<405> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1119 cl<404> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1120 cl<412> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1121 cl<413> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1122 cl<415> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1123 cl<414> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1124 cl<410> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1125 cl<411> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1126 cl<409> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1127 cl<408> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1128 cl<392> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1129 cl<393> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1130 cl<395> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1131 cl<394> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1132 cl<398> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1133 cl<399> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1134 cl<397> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1135 cl<388> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1136 cl<389> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1137 cl<391> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1138 cl<396> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1139 cl<390> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1140 cl<386> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1141 cl<387> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1142 cl<419> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1143 cl<418> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1144 cl<422> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1145 cl<428> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1146 cl<423> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1147 cl<421> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1148 cl<420> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1149 cl<429> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1150 cl<431> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1151 cl<430> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1152 cl<426> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1153 cl<427> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1154 cl<425> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1155 cl<424> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1156 cl<440> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1157 cl<441> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1158 cl<443> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1159 cl<442> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1160 cl<446> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1161 cl<447> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1162 cl<445> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1163 cl<444> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1164 cl<436> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1165 cl<437> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1166 cl<439> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1167 cl<438> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1168 cl<434> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1169 cl<435> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1170 cl<433> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1171 cl<432> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1172 cl<416> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1173 cl<417> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1174 cl<481> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1175 cl<480> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1176 cl<496> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1177 cl<497> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1178 cl<499> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1179 cl<498> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1180 cl<502> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1181 cl<503> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1182 cl<501> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1183 cl<500> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1184 cl<508> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1185 cl<509> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1186 cl<511> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1187 cl<510> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1188 cl<506> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1189 cl<507> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1190 cl<505> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1191 cl<504> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1192 cl<488> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1193 cl<489> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1194 cl<491> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1195 cl<490> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1196 cl<494> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1197 cl<495> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1198 cl<493> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1199 cl<484> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1200 cl<485> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1201 cl<487> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1202 cl<492> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1203 cl<486> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1204 cl<482> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1205 cl<483> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1206 cl<451> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1207 cl<450> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1208 cl<454> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1209 cl<460> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1210 cl<455> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1211 cl<453> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1212 cl<452> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1213 cl<461> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1214 cl<463> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1215 cl<462> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1216 cl<458> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1217 cl<459> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1218 cl<457> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1219 cl<456> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1220 cl<472> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1221 cl<473> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1222 cl<475> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1223 cl<474> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1224 cl<478> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1225 cl<479> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1226 cl<477> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1227 cl<476> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1228 cl<468> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1229 cl<469> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1230 cl<471> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1231 cl<470> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1232 cl<466> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1233 cl<467> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1234 cl<465> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1235 cl<464> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1236 cl<448> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1237 cl<449> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1238 cl<321> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1239 cl<320> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1240 cl<336> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1241 cl<337> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1242 cl<339> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1243 cl<338> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1244 cl<342> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1245 cl<343> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1246 cl<341> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1247 cl<340> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1248 cl<348> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1249 cl<349> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1250 cl<351> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1251 cl<350> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1252 cl<346> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1253 cl<347> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1254 cl<345> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1255 cl<344> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1256 cl<328> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1257 cl<329> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1258 cl<331> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1259 cl<330> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1260 cl<334> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1261 cl<335> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1262 cl<333> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1263 cl<324> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1264 cl<325> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1265 cl<327> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1266 cl<332> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1267 cl<326> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1268 cl<322> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1269 cl<323> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1270 cl<355> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1271 cl<354> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1272 cl<358> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1273 cl<364> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1274 cl<359> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1275 cl<357> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1276 cl<356> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1277 cl<365> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1278 cl<367> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1279 cl<366> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1280 cl<362> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1281 cl<363> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1282 cl<361> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1283 cl<360> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1284 cl<376> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1285 cl<377> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1286 cl<379> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1287 cl<378> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1288 cl<382> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1289 cl<383> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1290 cl<381> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1291 cl<380> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1292 cl<372> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1293 cl<373> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1294 cl<375> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1295 cl<374> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1296 cl<370> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1297 cl<371> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1298 cl<369> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1299 cl<368> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1300 cl<352> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1301 cl<353> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1302 cl<289> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1303 cl<288> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1304 cl<304> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1305 cl<305> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1306 cl<307> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1307 cl<306> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1308 cl<310> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1309 cl<311> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1310 cl<309> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1311 cl<308> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1312 cl<316> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1313 cl<317> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1314 cl<319> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1315 cl<318> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1316 cl<314> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1317 cl<315> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1318 cl<313> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1319 cl<312> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1320 cl<296> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1321 cl<297> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1322 cl<299> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1323 cl<298> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1324 cl<302> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1325 cl<303> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1326 cl<301> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1327 cl<292> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1328 cl<293> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1329 cl<295> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1330 cl<300> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1331 cl<294> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1332 cl<290> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1333 cl<291> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1334 cl<259> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1335 cl<258> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1336 cl<262> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1337 cl<268> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1338 cl<263> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1339 cl<261> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1340 cl<260> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1341 cl<269> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1342 cl<271> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1343 cl<270> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1344 cl<266> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1345 cl<267> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1346 cl<265> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1347 cl<264> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1348 cl<280> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1349 cl<281> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1350 cl<283> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1351 cl<282> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1352 cl<286> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1353 cl<287> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1354 cl<285> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1355 cl<284> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1356 cl<276> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1357 cl<277> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1358 cl<279> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1359 cl<278> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1360 cl<274> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1361 cl<275> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1362 cl<273> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1363 cl<272> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1364 cl<256> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI1365 cl<257> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI886 cl<35> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI854 cl<0> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
XI855 cl<1> net9403 net9404 l_sel n_ena p_ena pre r_sel wl<511> wl<510>
+wl<509> wl<508> wl<507> wl<506> wl<505> wl<504> wl<503> wl<502> wl<501>
+wl<500> wl<499> wl<498> wl<497> wl<496> wl<495> wl<494> wl<493> wl<492>
+wl<491> wl<490> wl<489> wl<488> wl<487> wl<486> wl<485> wl<484> wl<483>
+wl<482> wl<481> wl<480> wl<479> wl<478> wl<477> wl<476> wl<475> wl<474>
+wl<473> wl<472> wl<471> wl<470> wl<469> wl<468> wl<467> wl<466> wl<465>
+wl<464> wl<463> wl<462> wl<461> wl<460> wl<459> wl<458> wl<457> wl<456>
+wl<455> wl<454> wl<453> wl<452> wl<451> wl<450> wl<449> wl<448> wl<447>
+wl<446> wl<445> wl<444> wl<443> wl<442> wl<441> wl<440> wl<439> wl<438>
+wl<437> wl<436> wl<435> wl<434> wl<433> wl<432> wl<431> wl<430> wl<429>
+wl<428> wl<427> wl<426> wl<425> wl<424> wl<423> wl<422> wl<421> wl<420>
+wl<419> wl<418> wl<417> wl<416> wl<415> wl<414> wl<413> wl<412> wl<411>
+wl<410> wl<409> wl<408> wl<407> wl<406> wl<405> wl<404> wl<403> wl<402>
+wl<401> wl<400> wl<399> wl<398> wl<397> wl<396> wl<395> wl<394> wl<393>
+wl<392> wl<391> wl<390> wl<389> wl<388> wl<387> wl<386> wl<385> wl<384>
+wl<383> wl<382> wl<381> wl<380> wl<379> wl<378> wl<377> wl<376> wl<375>
+wl<374> wl<373> wl<372> wl<371> wl<370> wl<369> wl<368> wl<367> wl<366>
+wl<365> wl<364> wl<363> wl<362> wl<361> wl<360> wl<359> wl<358> wl<357>
+wl<356> wl<355> wl<354> wl<353> wl<352> wl<351> wl<350> wl<349> wl<348>
+wl<347> wl<346> wl<345> wl<344> wl<343> wl<342> wl<341> wl<340> wl<339>
+wl<338> wl<337> wl<336> wl<335> wl<334> wl<333> wl<332> wl<331> wl<330>
+wl<329> wl<328> wl<327> wl<326> wl<325> wl<324> wl<323> wl<322> wl<321>
+wl<320> wl<319> wl<318> wl<317> wl<316> wl<315> wl<314> wl<313> wl<312>
+wl<311> wl<310> wl<309> wl<308> wl<307> wl<306> wl<305> wl<304> wl<303>
+wl<302> wl<301> wl<300> wl<299> wl<298> wl<297> wl<296> wl<295> wl<294>
+wl<293> wl<292> wl<291> wl<290> wl<289> wl<288> wl<287> wl<286> wl<285>
+wl<284> wl<283> wl<282> wl<281> wl<280> wl<279> wl<278> wl<277> wl<276>
+wl<275> wl<274> wl<273> wl<272> wl<271> wl<270> wl<269> wl<268> wl<267>
+wl<266> wl<265> wl<264> wl<263> wl<262> wl<261> wl<260> wl<259> wl<258>
+wl<257> wl<256> wl<255> wl<254> wl<253> wl<252> wl<251> wl<250> wl<249>
+wl<248> wl<247> wl<246> wl<245> wl<244> wl<243> wl<242> wl<241> wl<240>
+wl<239> wl<238> wl<237> wl<236> wl<235> wl<234> wl<233> wl<232> wl<231>
+wl<230> wl<229> wl<228> wl<227> wl<226> wl<225> wl<224> wl<223> wl<222>
+wl<221> wl<220> wl<219> wl<218> wl<217> wl<216> wl<215> wl<214> wl<213>
+wl<212> wl<211> wl<210> wl<209> wl<208> wl<207> wl<206> wl<205> wl<204>
+wl<203> wl<202> wl<201> wl<200> wl<199> wl<198> wl<197> wl<196> wl<195>
+wl<194> wl<193> wl<192> wl<191> wl<190> wl<189> wl<188> wl<187> wl<186>
+wl<185> wl<184> wl<183> wl<182> wl<181> wl<180> wl<179> wl<178> wl<177>
+wl<176> wl<175> wl<174> wl<173> wl<172> wl<171> wl<170> wl<169> wl<168>
+wl<167> wl<166> wl<165> wl<164> wl<163> wl<162> wl<161> wl<160> wl<159>
+wl<158> wl<157> wl<156> wl<155> wl<154> wl<153> wl<152> wl<151> wl<150>
+wl<149> wl<148> wl<147> wl<146> wl<145> wl<144> wl<143> wl<142> wl<141>
+wl<140> wl<139> wl<138> wl<137> wl<136> wl<135> wl<134> wl<133> wl<132>
+wl<131> wl<130> wl<129> wl<128> wl<127> wl<126> wl<125> wl<124> wl<123>
+wl<122> wl<121> wl<120> wl<119> wl<118> wl<117> wl<116> wl<115> wl<114>
+wl<113> wl<112> wl<111> wl<110> wl<109> wl<108> wl<107> wl<106> wl<105>
+wl<104> wl<103> wl<102> wl<101> wl<100> wl<99> wl<98> wl<97> wl<96> wl<95>
+wl<94> wl<93> wl<92> wl<91> wl<90> wl<89> wl<88> wl<87> wl<86> wl<85> wl<84>
+wl<83> wl<82> wl<81> wl<80> wl<79> wl<78> wl<77> wl<76> wl<75> wl<74> wl<73>
+wl<72> wl<71> wl<70> wl<69> wl<68> wl<67> wl<66> wl<65> wl<64> wl<63> wl<62>
+wl<61> wl<60> wl<59> wl<58> wl<57> wl<56> wl<55> wl<54> wl<53> wl<52> wl<51>
+wl<50> wl<49> wl<48> wl<47> wl<46> wl<45> wl<44> wl<43> wl<42> wl<41> wl<40>
+wl<39> wl<38> wl<37> wl<36> wl<35> wl<34> wl<33> wl<32> wl<31> wl<30> wl<29>
+wl<28> wl<27> wl<26> wl<25> wl<24> wl<23> wl<22> wl<21> wl<20> wl<19> wl<18>
+wl<17> wl<16> wl<15> wl<14> wl<13> wl<12> wl<11> wl<10> wl<9> wl<8> wl<7>
+wl<6> wl<5> wl<4> wl<3> wl<2> wl<1> wl<0>   array512x1
.ENDS

************************************************************************
* Library Name: Lassen_DRAMB
* Cell Name: decoder6_64
* View Name: schematic
************************************************************************

.SUBCKT decoder6_64 A<5> A<4> A<3> A<2> A<1> A<0> ENA X<63> X<62> X<61> X<60>
+X<59> X<58> X<57> X<56> X<55> X<54> X<53> X<52> X<51> X<50> X<49> X<48> X<47>
+X<46> X<45> X<44> X<43> X<42> X<41> X<40> X<39> X<38> X<37> X<36> X<35> X<34>
+X<33> X<32> X<31> X<30> X<29> X<28> X<27> X<26> X<25> X<24> X<23> X<22> X<21>
+X<20> X<19> X<18> X<17> X<16> X<15> X<14> X<13> X<12> X<11> X<10> X<9> X<8>
+X<7> X<6> X<5> X<4> X<3> X<2> X<1> X<0>
XI95 A<5> A<4> ENA en<3> en<2> en<1> en<0>   decoder2_4
XI97 A<3> A<2> A<1> A<0> en<2> X<47> X<46> X<45> X<44> X<43> X<42> X<41> X<40>
+X<39> X<38> X<37> X<36> X<35> X<34> X<33> X<32>   decoder4_16
XI98 A<3> A<2> A<1> A<0> en<3> X<63> X<62> X<61> X<60> X<59> X<58> X<57> X<56>
+X<55> X<54> X<53> X<52> X<51> X<50> X<49> X<48>   decoder4_16
XI94 A<3> A<2> A<1> A<0> en<0> X<15> X<14> X<13> X<12> X<11> X<10> X<9> X<8>
+X<7> X<6> X<5> X<4> X<3> X<2> X<1> X<0>   decoder4_16
XI96 A<3> A<2> A<1> A<0> en<1> X<31> X<30> X<29> X<28> X<27> X<26> X<25> X<24>
+X<23> X<22> X<21> X<20> X<19> X<18> X<17> X<16>   decoder4_16
.ENDS

************************************************************************
* Library Name: Lassen_DRAMB
* Cell Name: bank16mx1n
* View Name: schematic
************************************************************************

.SUBCKT bank16mx1n a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14>
+a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> ena
+i_o w_
XI66 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<22> i_o w_   block512x512n
XI65 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<6> i_o w_   block512x512n
XI64 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<23> i_o w_   block512x512n
XI63 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<7> i_o w_   block512x512n
XI62 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<8> i_o w_   block512x512n
XI61 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<25> i_o w_   block512x512n
XI59 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<27> i_o w_   block512x512n
XI58 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<24> i_o w_   block512x512n
XI57 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<20> i_o w_   block512x512n
XI56 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<21> i_o w_   block512x512n
XI55 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<26> i_o w_   block512x512n
XI54 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<4> i_o w_   block512x512n
XI53 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<11> i_o w_   block512x512n
XI52 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<5> i_o w_   block512x512n
XI49 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<10> i_o w_   block512x512n
XI35 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<39> i_o w_   block512x512n
XI36 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<40> i_o w_   block512x512n
XI41 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<52> i_o w_   block512x512n
XI32 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<54> i_o w_   block512x512n
XI47 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<41> i_o w_   block512x512n
XI51 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<9> i_o w_   block512x512n
XI38 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<59> i_o w_   block512x512n
XI48 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<42> i_o w_   block512x512n
XI18 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<33> i_o w_   block512x512n
XI21 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<62> i_o w_   block512x512n
XI20 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<32> i_o w_   block512x512n
XI42 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<53> i_o w_   block512x512n
XI22 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<49> i_o w_   block512x512n
XI28 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<35> i_o w_   block512x512n
XI31 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<50> i_o w_   block512x512n
XI27 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<44> i_o w_   block512x512n
XI25 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<63> i_o w_   block512x512n
XI30 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<34> i_o w_   block512x512n
XI19 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<47> i_o w_   block512x512n
XI26 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<61> i_o w_   block512x512n
XI24 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<60> i_o w_   block512x512n
XI34 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<55> i_o w_   block512x512n
XI23 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<48> i_o w_   block512x512n
XI17 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<45> i_o w_   block512x512n
XI3 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<14> i_o w_   block512x512n
XI5 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<13> i_o w_   block512x512n
XI2 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<1> i_o w_   block512x512n
XI1 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<15> i_o w_   block512x512n
XI0 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<0> i_o w_   block512x512n
XI11 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<30> i_o w_   block512x512n
XI10 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<17> i_o w_   block512x512n
XI8 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<16> i_o w_   block512x512n
XI15 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<28> i_o w_   block512x512n
XI9 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<31> i_o w_   block512x512n
XI13 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<29> i_o w_   block512x512n
XI7 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<12> i_o w_   block512x512n
XI6 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<3> i_o w_   block512x512n
XI14 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<19> i_o w_   block512x512n
XI4 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<2> i_o w_   block512x512n
XI12 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<18> i_o w_   block512x512n
XI39 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<56> i_o w_   block512x512n
XI16 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<46> i_o w_   block512x512n
XI37 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<57> i_o w_   block512x512n
XI29 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<51> i_o w_   block512x512n
XI43 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<58> i_o w_   block512x512n
XI45 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<43> i_o w_   block512x512n
XI46 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<37> i_o w_   block512x512n
XI33 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<38> i_o w_   block512x512n
XI44 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> en<36> i_o w_   block512x512n
XI68 a<23> a<22> a<21> a<20> a<19> a<18> ena en<63> en<62> en<61> en<60>
+en<59> en<58> en<57> en<56> en<55> en<54> en<53> en<52> en<51> en<50> en<49>
+en<48> en<47> en<46> en<45> en<44> en<43> en<42> en<41> en<40> en<39> en<38>
+en<37> en<36> en<35> en<34> en<33> en<32> en<31> en<30> en<29> en<28> en<27>
+en<26> en<25> en<24> en<23> en<22> en<21> en<20> en<19> en<18> en<17> en<16>
+en<15> en<14> en<13> en<12> en<11> en<10> en<9> en<8> en<7> en<6> en<5> en<4>
+en<3> en<2> en<1> en<0>   decoder6_64
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: atd18
* View Name: schematic
************************************************************************

.SUBCKT atd18 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7>
+a<6> a<5> a<4> a<3> a<2> a<1> a<0> w_ y
XI103 net99 net97 net189 net163   nor3 Lp=0.35u Wp=7u Ln=0.35u Wn=3.5u
XI74 net157 net152 net147 net142 net163 net137   nand5 Lp=0.35u Wp=4u Ln=0.35u
+Wn=7u
XI96 net169 net165 net171 net167 net142   nor4 Lp=0.35u Wp=7u Ln=0.35u Wn=3.5u
XI93 net181 net183 net187 net185 net152   nor4 Lp=0.35u Wp=7u Ln=0.35u Wn=3.5u
XI92 net193 net195 net197 net191 net157   nor4 Lp=0.35u Wp=7u Ln=0.35u Wn=3.5u
XI94 net175 net179 net173 net177 net147   nor4 Lp=0.35u Wp=7u Ln=0.35u Wn=3.5u
XI75 net137 net159   inv Ln=0.35u Wn=8u M=3 Lp=0.35u Wp=16u
XI81 net159 y   inv Ln=0.35u Wn=8u M=9 Lp=0.35u Wp=16u
XI101 a<16> net99   atd1
XI102 a<17> net97   atd1
XI97 a<14> net171   atd1
XI98 a<12> net169   atd1
XI71 a<3> net191   atd1
XI99 a<15> net167   atd1
XI79 w_ net189   atd1
XI91 a<10> net173   atd1
XI68 a<0> net193   atd1
XI83 a<4> net181   atd1
XI84 a<5> net183   atd1
XI82 a<7> net185   atd1
XI88 a<8> net175   atd1
XI85 a<6> net187   atd1
XI100 a<13> net165   atd1
XI69 a<1> net195   atd1
XI70 a<2> net197   atd1
XI90 a<11> net177   atd1
XI89 a<9> net179   atd1
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: dff1
* View Name: schematic
************************************************************************

.SUBCKT dff1 clk d q
XI71 net46 net30   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI80 clk ck_   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI81 ck_ ck   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI75 net30 net42   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI77 q net38   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI76 net34 q   inv Ln=0.35u Wn=7u M=1 Lp=0.35u Wp=14u
XI73 d net46 ck_ ck   ctg Lp=0.35u Wp=3.5u Ln=0.35u Wn=3.5u
XI74 net46 net42 ck ck_   ctg Lp=0.35u Wp=3.5u Ln=0.35u Wn=3.5u
XI78 net34 net38 ck_ ck   ctg Lp=0.35u Wp=3.5u Ln=0.35u Wn=3.5u
XI79 net30 net34 ck ck_   ctg Lp=0.35u Wp=3.5u Ln=0.35u Wn=3.5u
.ENDS

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: level_shift1
* View Name: schematic
************************************************************************

.SUBCKT level_shift1 IN OUT VDD VSS
M1 tn1 OUT VDD VDD PMOS W=3.5u L=350.00n M=1
M2 OUT tn1 VDD VDD PMOS W=3.5u L=350.00n M=1
M3 tn1 IN VSS VSS NMOS W=1.4u L=350.00n M=1
M4 OUT INB VSS VSS NMOS W=1.4u L=350.00n M=1
XIV1 IN INB inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
.ENDS level_shift1

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: level_shift2
* View Name: schematic
************************************************************************

.SUBCKT level_shift2 IN OUT VDD VSS
M1 tn1 OUT VDD VDD PMOS W=3.5u L=350.00n M=1
M2 tn2 tn3 VDD VDD PMOS W=3.5u L=350.00n M=1
M3 tn3 IN tn1 VDD PMOS W=3.5u L=350.00n M=1
M4 OUT INB tn2 VDD PMOS W=3.5u L=350.00n M=1
M5 tn3 IN VSS VSS NMOS W=1.4u L=350.00n M=1
M6 OUT INB VSS VSS NMOS W=1.4u L=350.00n M=1
XIV1 IN INB inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
.ENDS level_shift2

************************************************************************
* Library Name: Lassen_DRAM
* Cell Name: level_shift3
* View Name: schematic
************************************************************************

.SUBCKT level_shift3 IN OUT VDD VBIASH VBIASL VSS
M1 tn1 tn2 VDD VDD PMOS W=3.5u L=350.00n M=1
M2 tn2 tn1 VDD VDD PMOS W=3.5u L=350.00n M=1
M3 tn3 VBIASH tn1 VDD PMOS W=3.5u L=350.00n M=1
M4 OUT VBIASH tn2 VDD PMOS W=3.5u L=350.00n M=1
M5 tn3 VBIASL tn5 VSS NMOS W=1.4u L=350.00n M=1
M6 OUT VBIASL tn6 VSS NMOS W=1.4u L=350.00n M=1
M7 tn5 INB VSS VSS NMOS W=1.4u L=350.00n M=1
M8 tn6 IN VSS VSS NMOS W=1.4u L=350.00n M=1
XIV1 IN INB inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
.ENDS level_shift3

************************************************************************
* Library Name: Lassen_DRAMB
* Cell Name: dram1gbn
* View Name: schematic
************************************************************************

.SUBCKT dram1gbn a<29> a<28> a<27> a<26> a<25> a<24> a<23> a<22> a<21> a<20>
+a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7>
+a<6> a<5> a<4> a<3> a<2> a<1> a<0> d ena q w_
XI66 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<22> 0 net230
+  bank16mx1n
XI65 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<6> 0 net230
+  bank16mx1n
XI64 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<23> 0 net230
+  bank16mx1n
XI63 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<7> 0 net230
+  bank16mx1n
XI62 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<8> 0 net230
+  bank16mx1n
XI61 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<25> 0 net230
+  bank16mx1n
XI59 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<27> 0 net230
+  bank16mx1n
XI58 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<24> 0 net230
+  bank16mx1n
***XI57 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<20> 0 net230
***+  bank16mx1n
***XI56 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<21> 0 net230
***+  bank16mx1n
***XI55 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<26> 0 net230
***+  bank16mx1n
***XI54 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<4> 0 net230
***+  bank16mx1n
***XI53 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<11> 0 net230
***+  bank16mx1n
***XI52 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<5> 0 net230
***+  bank16mx1n
***XI49 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<10> 0 net230
***+  bank16mx1n
***XI35 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<39> 0 net230
***+  bank16mx1n
***XI36 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<40> 0 net230
***+  bank16mx1n
***XI41 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<52> 0 net230
***+  bank16mx1n
***XI32 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<54> 0 net230
***+  bank16mx1n
***XI47 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<41> 0 net230
***+  bank16mx1n
***XI51 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<9> 0 net230
***+  bank16mx1n
***XI38 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<59> 0 net230
***+  bank16mx1n
***XI48 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<42> 0 net230
***+  bank16mx1n
***XI18 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<33> 0 net230
***+  bank16mx1n
***XI21 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<62> 0 net230
***+  bank16mx1n
***XI20 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<32> 0 net230
***+  bank16mx1n
***XI42 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<53> 0 net230
***+  bank16mx1n
***XI22 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<49> 0 net230
***+  bank16mx1n
***XI28 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<35> 0 net230
***+  bank16mx1n
***XI31 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<50> 0 net230
***+  bank16mx1n
***XI27 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<44> 0 net230
***+  bank16mx1n
***XI25 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<63> 0 net230
***+  bank16mx1n
***XI30 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<34> 0 net230
***+  bank16mx1n
***XI19 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<47> 0 net230
***+  bank16mx1n
***XI26 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<61> 0 net230
***+  bank16mx1n
***XI24 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<60> 0 net230
***+  bank16mx1n
***XI34 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<55> 0 net230
***+  bank16mx1n
***XI23 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<48> 0 net230
***+  bank16mx1n
***XI17 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<45> 0 net230
***+  bank16mx1n
***XI3 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<14> 0 net230
***+  bank16mx1n
***XI5 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<13> 0 net230
***+  bank16mx1n
***XI2 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<1> 0 net230
***+  bank16mx1n
***XI1 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<15> 0 net230
***+  bank16mx1n
***XI0 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<0> io_x net230
***+  bank16mx1n
***XI11 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<30> 0 net230
***+  bank16mx1n
***XI10 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<17> 0 net230
***+  bank16mx1n
***XI8 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<16> 0 net230
***+  bank16mx1n
***XI15 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<28> 0 net230
***+  bank16mx1n
***XI9 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<31> 0 net230
***+  bank16mx1n
***XI13 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<29> 0 net230
***+  bank16mx1n
***XI7 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<12> 0 net230
***+  bank16mx1n
***XI6 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<3> 0 net230
***+  bank16mx1n
***XI14 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<19> 0 net230
***+  bank16mx1n
***XI4 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<2> 0 net230
***+  bank16mx1n
***XI12 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<18> 0 net230
***+  bank16mx1n
***XI39 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<56> 0 net230
***+  bank16mx1n
***XI16 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<46> 0 net230
***+  bank16mx1n
***XI37 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<57> 0 net230
***+  bank16mx1n
***XI29 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<51> 0 net230
***+  bank16mx1n
***XI43 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<58> 0 net230
***+  bank16mx1n
***XI45 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<43> 0 net230
***+  bank16mx1n
***XI46 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<37> 0 net230
***+  bank16mx1n
***XI33 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<38> 0 net230
***+  bank16mx1n
***XI44 a<23> a<22> a<21> a<20> a<19> a<18> a<17> a<16> a<15> a<14> a<13> a<12>
***+a<11> a<10> a<9> a<8> a<7> a<6> a<5> a<4> a<3> a<2> a<1> a<0> en<36> 0 net230
***+  bank16mx1n
XI73 a<17> a<16> a<15> a<14> a<13> a<12> a<11> a<10> a<9> a<8> a<7> a<6> a<5>
+a<4> a<3> a<2> a<1> a<0> net230 net474   atd18
XI160 net476 net493   inv Ln=0.35u Wn=20u M=2 Lp=0.35u Wp=40u
XI310 w_ net480   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI309 net480 net230   inv Ln=0.35u Wn=20u M=2 Lp=0.35u Wp=40u
XI83 d net476   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI221 net491 net485   inv Ln=0.35u Wn=7u M=6 Lp=0.35u Wp=14u
XI159 net230 net487   inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u
XI222 net485 q   inv Ln=0.35u Wn=7u M=12 Lp=0.35u Wp=14u
XI223 net496 net491   inv Ln=0.35u Wn=7u M=2 Lp=0.35u Wp=14u
XI161 io_x net493 net487 net230   ctg Lp=0.35u Wp=3.5u Ln=0.35u Wn=3.5u
XI74 net500 io_x  net496   dff1
XI72 net501 net500 net503   sen_ena
XI71 net474 net503   xvald
XI68 a<29> a<28> a<27> a<26> a<25> a<24> ena en<63> en<62> en<61> en<60>
+en<59> en<58> en<57> en<56> en<55> en<54> en<53> en<52> en<51> en<50> en<49>
+en<48> en<47> en<46> en<45> en<44> en<43> en<42> en<41> en<40> en<39> en<38>
+en<37> en<36> en<35> en<34> en<33> en<32> en<31> en<30> en<29> en<28> en<27>
+en<26> en<25> en<24> en<23> en<22> en<21> en<20> en<19> en<18> en<17> en<16>
+en<15> en<14> en<13> en<12> en<11> en<10> en<9> en<8> en<7> en<6> en<5> en<4>
+en<3> en<2> en<1> en<0>   decoder6_64
.ENDS