.SUBCKT rl_sel a pre sel xvld
XI41 pre pre_out  inv Ln=0.35u Wn=4u M=1 Lp=0.35u Wp=8u

MM14 net28 xvld gnd! vbb! NMOS W=8u L=0.35u M=1
MM13 Y A net28 vbb! NMOS W=8u L=0.35u M=1
MM12 Y A vddh2! vddh2! PMOS W=4u L=0.35u M=1.0
MM11 Y xvld vddh2! vddh2! PMOS W=4u L=0.35u M=1.0

MM15 i1 Y gnd! vbb! NMOS W=14u L=350.00n M=1
MM6  i1 Y vddh2! vddh2! PMOS W=28u L=350.00n M=1.0
MM16 i2 i1 gnd! vbb! NMOS W=14u L=350.00n M=1
MM7  i2 i1 vddh2! vddh2! PMOS W=28u L=350.00n M=1.0
MM17 sel i2 gnd! vbb! NMOS W=14u L=350.00n M=1
MM8  sel i2 vddh2! vddh2! PMOS W=28u L=350.00n M=1.0
.ENDS
